* NGSPICE file created from CM.ext - technology: gf180mcuD

.subckt CM VREF VB VSS VCOPY
X0 VCOPY VREF VSS VSUBS nfet_03v3 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=1.41u
X1 a_n2186_n1122# a_n2186_n1122# a_n2186_n1122# VSUBS nfet_03v3 ad=1.856p pd=7.56u as=30.7232p ps=0.15968m w=3.2u l=1.41u
X2 VCOPY VREF VSS VSUBS nfet_03v3 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=1.41u
X3 VREF VREF VSS VSUBS nfet_03v3 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=1.41u
X4 a_n2186_n1122# a_n2186_n1122# a_n2186_n1122# VSUBS nfet_03v3 ad=1.856p pd=7.56u as=0 ps=0 w=3.2u l=1.41u
X5 VREF VREF VSS VSUBS nfet_03v3 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=1.41u
C0 VCOPY VREF 0.44525f
C1 VCOPY VSS 2.51605f
C2 VCOPY a_n2186_n1122# 1.23099f
C3 VB VREF 0
C4 VB VSS 0.00158f
C5 VB a_n2186_n1122# 0.04115f
C6 VREF VSS 4.6056f
C7 a_n2186_n1122# VREF 1.34245f
C8 a_n2186_n1122# VSS 0.52287f
C9 VCOPY VB 0.00304f
C10 VB VSUBS 0.02607f
C11 VCOPY VSUBS 0.83945f
C12 VSS VSUBS 1.63231f
C13 VREF VSUBS 4.7845f
C14 a_n2186_n1122# VSUBS 7.80005f
.ends

