* Extracted by KLayout with GF180MCU LVS runset on : 24/09/2025 18:46

.SUBCKT TOP
M$1 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$2 \$247 \$247 \$269 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$3 \$252 \$247 \$251 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$4 \$254 \$247 \$253 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$5 \$256 \$247 \$255 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$6 VIN_OUT \$247 \$257 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$7 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$8 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$9 \$269 \$269 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$10 \$251 \$269 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$11 \$253 \$269 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$12 \$255 \$269 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$13 \$257 \$269 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$14 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$15 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$16 \$351 \$351 \$360 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$17 \$351 \$351 \$360 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$18 \$351 \$351 \$360 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$19 \$351 \$351 \$360 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$20 \$351 \$351 \$360 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$21 \$351 \$351 \$360 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$22 \$351 \$351 \$360 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$23 \$351 \$351 \$360 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$24 \$351 \$351 \$360 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$25 \$351 \$351 \$360 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$26 \$362 \$351 \$361 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$27 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$28 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$29 \$352 \$352 \$363 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$30 \$352 \$352 \$363 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$31 \$352 \$352 \$363 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$32 \$352 \$352 \$363 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$33 \$352 \$352 \$363 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$34 \$352 \$352 \$363 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$35 \$352 \$352 \$363 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$36 \$352 \$352 \$363 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$37 \$352 \$352 \$363 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$38 \$352 \$352 \$363 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$39 \$320 \$352 \$364 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$40 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$41 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$42 \$269 \$313 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$43 \$269 \$313 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$44 \$269 \$313 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$45 \$269 \$313 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$46 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$47 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$48 \$360 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$49 \$360 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$50 \$360 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$51 \$360 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$52 \$360 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$53 \$360 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$54 \$360 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$55 \$360 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$56 \$360 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$57 \$360 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$58 \$361 \$360 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$59 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$60 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$61 \$363 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$62 \$363 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$63 \$363 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$64 \$363 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$65 \$363 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$66 \$363 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$67 \$363 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$68 \$363 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$69 \$363 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$70 \$363 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$71 \$364 \$363 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$72 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$73 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$74 \$360 \$313 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$75 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$76 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$77 \$363 \$313 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$78 VDD VDD VDD VDD pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P PS=21.16U PD=21.16U
M$79 \$204 \$169 \$203 \$210 pfet_05v0 L=0.5U W=0.9U AS=0.396P AD=0.396P
+ PS=2.68U PD=2.68U
M$80 \$204 \$168 \$168 \$217 pfet_05v0 L=0.5U W=0.9U AS=0.396P AD=0.396P
+ PS=2.68U PD=2.68U
M$81 VSS VSS VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.64P AD=4.64P PS=17.16U
+ PD=17.16U
M$82 \$373 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$83 \$373 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$84 \$373 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$85 \$373 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$86 \$373 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$87 \$373 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$88 \$373 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$89 \$373 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$90 \$373 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$91 \$373 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$92 \$382 \$373 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$93 VSS VSS VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.64P AD=4.64P PS=17.16U
+ PD=17.16U
M$94 VSS VSS VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.64P AD=4.64P PS=17.16U
+ PD=17.16U
M$95 \$362 \$362 \$373 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$96 \$362 \$362 \$373 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$97 \$362 \$362 \$373 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$98 \$362 \$362 \$373 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$99 \$362 \$362 \$373 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$100 \$362 \$362 \$373 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$101 \$362 \$362 \$373 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$102 \$362 \$362 \$373 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$103 \$362 \$362 \$373 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$104 \$362 \$362 \$373 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$105 \$352 \$362 \$382 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$106 VSS VSS VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.64P AD=4.64P PS=17.16U
+ PD=17.16U
M$107 \$75 \$169 \$169 gf180mcu_gnd nfet_05v0 L=0.6U W=0.66U AS=0.2904P
+ AD=0.2904P PS=2.2U PD=2.2U
M$108 \$75 \$168 \$213 gf180mcu_gnd nfet_05v0 L=0.6U W=0.66U AS=0.2904P
+ AD=0.2904P PS=2.2U PD=2.2U
M$109 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$110 \$252 \$252 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$111 VCM_OUT \$252 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$112 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$113 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$114 \$272 \$272 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$115 \$292 \$272 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$116 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$117 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$118 \$254 \$254 \$272 VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$119 BCM_OUT \$254 \$292 VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$120 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$121 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$122 CCM_OUT \$320 \$318 VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$123 \$320 \$318 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$124 CCM_OUT \$320 \$318 VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$125 \$320 \$318 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$126 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$127 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$128 \$353 \$256 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$129 \$318 \$256 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$130 \$353 \$256 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$131 \$318 \$256 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$132 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$133 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
M$134 \$320 \$353 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$135 \$256 \$320 \$353 VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$136 \$320 \$353 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$137 \$256 \$320 \$353 VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$138 VSS VSS VSS VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P PS=9.16U PD=9.16U
D$139 VSS \$74 diode_nd2ps_06v0 A=100P P=40U
D$140 VSS \$74 diode_nd2ps_06v0 A=100P P=40U
D$141 VSS \$74 diode_nd2ps_06v0 A=100P P=40U
D$142 VSS \$74 diode_nd2ps_06v0 A=100P P=40U
D$143 VSS \$225 diode_nd2ps_06v0 A=100P P=40U
D$144 VSS \$225 diode_nd2ps_06v0 A=100P P=40U
D$145 VSS \$225 diode_nd2ps_06v0 A=100P P=40U
D$146 VSS \$225 diode_nd2ps_06v0 A=100P P=40U
D$147 VSS \$322 diode_nd2ps_06v0 A=100P P=40U
D$148 VSS \$322 diode_nd2ps_06v0 A=100P P=40U
D$149 VSS \$322 diode_nd2ps_06v0 A=100P P=40U
D$150 VSS \$322 diode_nd2ps_06v0 A=100P P=40U
D$151 \$74 VDD diode_pd2nw_06v0 A=100P P=40U
D$152 \$74 VDD diode_pd2nw_06v0 A=100P P=40U
D$153 \$74 VDD diode_pd2nw_06v0 A=100P P=40U
D$154 \$74 VDD diode_pd2nw_06v0 A=100P P=40U
D$155 \$225 VDD diode_pd2nw_06v0 A=100P P=40U
D$156 \$225 VDD diode_pd2nw_06v0 A=100P P=40U
D$157 \$225 VDD diode_pd2nw_06v0 A=100P P=40U
D$158 \$225 VDD diode_pd2nw_06v0 A=100P P=40U
D$159 \$322 VDD diode_pd2nw_06v0 A=100P P=40U
D$160 \$322 VDD diode_pd2nw_06v0 A=100P P=40U
D$161 \$322 VDD diode_pd2nw_06v0 A=100P P=40U
D$162 \$322 VDD diode_pd2nw_06v0 A=100P P=40U
R$163 \$74 EN gf180mcu_gnd 87.5 ppolyf_u L=10U W=40U
R$164 \$225 VBIAS gf180mcu_gnd 87.5 ppolyf_u L=10U W=40U
R$165 \$322 VIN gf180mcu_gnd 87.5 ppolyf_u L=10U W=40U
.ENDS TOP
