| units: 0.5 tech: gf180mcuD format: MIT
x sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# VDD PD VDD s=15840,536 d=15840,536 l=100 w=180 x=514986 y=227349 pfet_05v0
x sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# TEXT$9_0/VSUBS sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# TEXT$9_0/VSUBS s=11616,440 d=11616,440 l=120 w=132 x=514986 y=227721 nfet_05v0
x sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# TEXT$9_0/VSUBS PU TEXT$9_0/VSUBS s=11616,440 d=11616,440 l=120 w=132 x=514985 y=226108 nfet_05v0
x sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# VDD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# VDD s=15840,536 d=15840,536 l=100 w=180 x=515005 y=226480 pfet_05v0
x io_secondary_5p0$1_0/ppolyf_u_9H3LNU_0/a_n224793_504155# EN m3_419992_265695# VDD s=816000,16204 d=816000,16204 l=2000 w=8000 x=510003 y=227557 ppolyf_u
x m3_419992_265695# TEXT$9_0/VSUBS l=0 w=0 x=503355 y=217079 diode_nd2ps_06v0
x m3_419992_265695# TEXT$9_0/VSUBS l=0 w=0 x=498891 y=217079 diode_nd2ps_06v0
x m3_419992_265695# TEXT$9_0/VSUBS l=0 w=0 x=501123 y=217079 diode_nd2ps_06v0
x m3_419992_265695# TEXT$9_0/VSUBS l=0 w=0 x=505587 y=217079 diode_nd2ps_06v0
x m3_419992_265695# VDD s=21168000,22704 l=0 w=0 x=498887 y=228335 diode_pd2nw_06v0
x m3_419992_265695# VDD s=21168000,22704 l=0 w=0 x=505535 y=228335 diode_pd2nw_06v0
x m3_419992_265695# VDD s=21168000,22704 l=0 w=0 x=501103 y=228335 diode_pd2nw_06v0
x m3_419992_265695# VDD s=21168000,22704 l=0 w=0 x=503319 y=228335 diode_pd2nw_06v0
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=387920 y=265903 pfet_03v3
x M_0/a_365708_259299# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=371358 y=262205 pfet_03v3
x M_0/a_365708_259299# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=367408 y=262205 pfet_03v3
x a_498947_268180# M_0/a_401941_244568# M_0/a_402461_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=402061 y=244568 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=366636 y=265903 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=400463 y=244568 pfet_03v3
x M_0/a_401151_244568# VDD M_0/a_404311_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=404431 y=249916 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=386304 y=262205 pfet_03v3
x a_499016_248165# M_0/a_373878_259299# M_0/a_374398_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=373998 y=259299 pfet_03v3
x M_0/a_386992_259299# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=388692 y=262205 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=396090 y=259299 pfet_03v3
x M_0/a_383940_262205# M_0/a_386992_259299# M_0/a_383940_262205# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=392642 y=259299 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=386304 y=265903 pfet_03v3
x M_0/a_401151_244568# VDD M_0/a_401151_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=401271 y=249916 pfet_03v3
x m4_400150_261569# M_0/a_409618_260539# M_0/a_404041_244568# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410208 y=260919 nfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=185600,3432 l=200 w=1600 x=376962 y=259699 nfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=411996 y=258781 nfet_03v3
x a_499016_248165# M_0/a_365708_259299# a_499016_248165# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=371358 y=259299 pfet_03v3
x M_0/a_409618_260539# TEXT$9_0/VSUBS m4_400150_261569# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=409618 y=260919 nfet_03v3
x a_499016_248165# M_0/a_365708_259299# a_499016_248165# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=367408 y=259299 pfet_03v3
x M_0/a_409498_256643# TEXT$9_0/VSUBS m4_400150_261569# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=411388 y=256643 nfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_377450_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=378750 y=259699 nfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=185600,3432 l=200 w=1600 x=376962 y=262205 nfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=411452 y=242557 nfet_03v3
x M_0/a_409618_260539# TEXT$9_0/VSUBS m4_400150_261569# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410798 y=260919 nfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_377450_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=378160 y=259699 nfet_03v3
x m3_419992_265695# VDD M_0/a_401151_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=401666 y=255368 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=386304 y=259299 pfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=185600,3432 l=200 w=1600 x=384348 y=259699 nfet_03v3
x M_0/a_365708_259299# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=372938 y=262205 pfet_03v3
x M_0/a_374398_259299# M_0/a_377450_262205# M_0/a_374398_259299# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=378750 y=262205 nfet_03v3
x m3_419992_265695# VDD M_0/a_401151_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=404036 y=255368 pfet_03v3
x M_0/a_383940_262205# M_0/a_386992_259299# M_0/a_383940_262205# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=388692 y=259299 pfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=409010 y=260919 nfet_03v3
x a_498947_268180# M_0/a_403521_244568# M_0/a_404041_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=403641 y=244568 pfet_03v3
x M_0/a_386992_259299# VDD M_0/a_395162_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=395282 y=262205 pfet_03v3
x M_0/a_386992_259299# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=393432 y=262205 pfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=409646 y=242557 nfet_03v3
x M_0/a_374398_259299# M_0/a_377450_262205# M_0/a_374398_259299# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=378160 y=262205 nfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_377450_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=382880 y=259699 nfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=185600,3432 l=200 w=1600 x=384348 y=262205 nfet_03v3
x M_0/a_365708_259299# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=372148 y=262205 pfet_03v3
x M_0/a_365708_259299# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=365828 y=262205 pfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_377450_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=382290 y=259699 nfet_03v3
x M_0/a_386992_259299# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=390272 y=262205 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=405239 y=249916 pfet_03v3
x M_0/a_374398_259299# M_0/a_377450_262205# M_0/a_374398_259299# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=382880 y=262205 nfet_03v3
x M_0/a_365708_259299# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=368988 y=262205 pfet_03v3
x M_0/a_401151_244568# VDD M_0/a_402731_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=402851 y=249916 pfet_03v3
x m3_419992_265695# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=365828 y=265903 pfet_03v3
x M_0/a_374398_259299# M_0/a_377450_262205# M_0/a_374398_259299# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=382290 y=262205 nfet_03v3
x a_499016_248165# M_0/a_365708_259299# a_499016_248165# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=372938 y=259299 pfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=411452 y=249599 nfet_03v3
x M_0/a_386992_259299# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=389482 y=262205 pfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=411452 y=251737 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=374806 y=262205 pfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=411996 y=256643 nfet_03v3
x M_0/a_404041_244568# TEXT$9_0/VSUBS M_0/a_409498_256643# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410208 y=258781 nfet_03v3
x M_0/a_383940_262205# M_0/a_395162_259299# m4_400150_261569# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=395282 y=259299 pfet_03v3
x M_0/a_383940_262205# M_0/a_386992_259299# M_0/a_383940_262205# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=393432 y=259299 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=365020 y=262205 pfet_03v3
x M_0/a_404041_244568# TEXT$9_0/VSUBS M_0/a_409618_260539# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=409618 y=258781 nfet_03v3
x M_0/a_401151_244568# VDD M_0/a_401941_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=402061 y=249916 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=404844 y=255368 pfet_03v3
x M_0/a_365708_259299# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=368198 y=262205 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=400463 y=249916 pfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=409646 y=249599 nfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=409646 y=251737 nfet_03v3
x a_499016_248165# M_0/a_365708_259299# a_499016_248165# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=372148 y=259299 pfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_377450_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=380520 y=259699 nfet_03v3
x a_499016_248165# M_0/a_365708_259299# a_499016_248165# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=365828 y=259299 pfet_03v3
x M_0/a_404041_244568# TEXT$9_0/VSUBS M_0/a_409618_260539# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410798 y=258781 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=365020 y=265903 pfet_03v3
x M_0/a_383940_262205# M_0/a_386992_259299# M_0/a_383940_262205# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=390272 y=259299 pfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_377450_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=379930 y=259699 nfet_03v3
x M_0/a_402461_244568# TEXT$9_0/VSUBS VCM_OUT TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410844 y=242557 nfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=409010 y=258781 nfet_03v3
x a_499016_248165# M_0/a_365708_259299# a_499016_248165# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=368988 y=259299 pfet_03v3
x m3_419992_265695# VDD M_0/a_401151_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=402456 y=255368 pfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_377450_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=379340 y=259699 nfet_03v3
x M_0/a_374398_259299# M_0/a_377450_262205# M_0/a_374398_259299# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=380520 y=262205 nfet_03v3
x M_0/a_402461_244568# TEXT$9_0/VSUBS M_0/a_402461_244568# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410254 y=242557 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=400858 y=255368 pfet_03v3
x M_0/a_383940_262205# M_0/a_386992_259299# M_0/a_383940_262205# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=389482 y=259299 pfet_03v3
x M_0/a_374398_259299# M_0/a_377450_262205# M_0/a_374398_259299# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=379930 y=262205 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=374806 y=259299 pfet_03v3
x m4_400150_261569# M_0/a_409618_260539# M_0/a_404041_244568# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=411388 y=260919 nfet_03v3
x M_0/a_386992_259299# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=391852 y=262205 pfet_03v3
x a_498947_268180# M_0/a_404311_244568# VIN_OUT VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=404431 y=244568 pfet_03v3
x M_0/a_386992_259299# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=394222 y=262205 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=365020 y=259299 pfet_03v3
x M_0/a_374398_259299# M_0/a_377450_262205# M_0/a_374398_259299# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=379340 y=262205 nfet_03v3
x M_0/a_386992_259299# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=387902 y=262205 pfet_03v3
x a_499016_248165# M_0/a_365708_259299# a_499016_248165# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=368198 y=259299 pfet_03v3
x M_0/a_365708_259299# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=370568 y=262205 pfet_03v3
x M_0/a_365708_259299# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=366618 y=262205 pfet_03v3
x a_498947_268180# M_0/a_401151_244568# a_498947_268180# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=401271 y=244568 pfet_03v3
x M_0/a_386992_259299# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=391062 y=262205 pfet_03v3
x M_0/a_401151_244568# VDD M_0/a_403521_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=403641 y=249916 pfet_03v3
x M_0/a_386992_259299# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=387112 y=262205 pfet_03v3
x M_0/a_365708_259299# VDD M_0/a_365708_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=369778 y=262205 pfet_03v3
x M_0/a_410134_251737# TEXT$9_0/VSUBS M_0/a_410724_251737# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410844 y=249599 nfet_03v3
x M_0/a_409498_256643# TEXT$9_0/VSUBS m4_400150_261569# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410208 y=256643 nfet_03v3
x M_0/a_403251_244568# M_0/a_410724_251737# BCM_OUT TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410844 y=251737 nfet_03v3
x m4_400150_261569# M_0/a_409498_256643# CCM_OUT TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=409618 y=256643 nfet_03v3
x m3_419992_265695# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=387112 y=265903 pfet_03v3
x M_0/a_383940_262205# M_0/a_386992_259299# M_0/a_383940_262205# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=391852 y=259299 pfet_03v3
x M_0/a_410134_251737# TEXT$9_0/VSUBS M_0/a_410134_251737# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410254 y=249599 nfet_03v3
x M_0/a_403251_244568# M_0/a_410134_251737# M_0/a_403251_244568# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410254 y=251737 nfet_03v3
x M_0/a_383940_262205# M_0/a_386992_259299# M_0/a_383940_262205# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=394222 y=259299 pfet_03v3
x M_0/a_383940_262205# M_0/a_386992_259299# M_0/a_383940_262205# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=387902 y=259299 pfet_03v3
x m4_400150_261569# M_0/a_409498_256643# CCM_OUT TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=410798 y=256643 nfet_03v3
x a_499016_248165# M_0/a_365708_259299# a_499016_248165# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=370568 y=259299 pfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=409010 y=256643 nfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_377450_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=381700 y=259699 nfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_377450_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=377570 y=259699 nfet_03v3
x a_499016_248165# M_0/a_365708_259299# a_499016_248165# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=366618 y=259299 pfet_03v3
x M_0/a_383940_262205# M_0/a_386992_259299# M_0/a_383940_262205# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=391062 y=259299 pfet_03v3
x TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS TEXT$9_0/VSUBS d=92800,1832 l=200 w=800 x=411996 y=260919 nfet_03v3
x M_0/a_383940_262205# M_0/a_386992_259299# M_0/a_383940_262205# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=387112 y=259299 pfet_03v3
x a_499016_248165# M_0/a_365708_259299# a_499016_248165# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=369778 y=259299 pfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_383620_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=383740 y=259699 nfet_03v3
x M_0/a_377450_262205# TEXT$9_0/VSUBS M_0/a_377450_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=381110 y=259699 nfet_03v3
x M_0/a_365708_259299# VDD M_0/a_373878_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=373998 y=262205 pfet_03v3
x M_0/a_374398_259299# M_0/a_377450_262205# M_0/a_374398_259299# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=377570 y=262205 nfet_03v3
x M_0/a_404041_244568# TEXT$9_0/VSUBS M_0/a_409498_256643# TEXT$9_0/VSUBS s=96000,1840 d=96000,1840 l=200 w=800 x=411388 y=258781 nfet_03v3
x m3_419992_265695# VDD M_0/a_401151_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=403246 y=255368 pfet_03v3
x M_0/a_374398_259299# M_0/a_377450_262205# M_0/a_374398_259299# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=381700 y=262205 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=405239 y=244568 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=396090 y=262205 pfet_03v3
x a_498947_268180# M_0/a_402731_244568# M_0/a_403251_244568# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=402851 y=244568 pfet_03v3
x M_0/a_386992_259299# VDD M_0/a_386992_259299# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=392642 y=262205 pfet_03v3
x M_0/a_374398_259299# M_0/a_383620_262205# M_0/a_383940_262205# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=383740 y=262205 nfet_03v3
x M_0/a_374398_259299# M_0/a_377450_262205# M_0/a_374398_259299# TEXT$9_0/VSUBS s=192000,3440 d=192000,3440 l=200 w=1600 x=381110 y=262205 nfet_03v3
x a_498947_268180# VDD s=21168000,22704 l=0 w=0 x=505595 y=268180 diode_pd2nw_06v0
x a_498947_268180# VDD s=21168000,22704 l=0 w=0 x=501163 y=268180 diode_pd2nw_06v0
x a_499016_248165# TEXT$9_0/VSUBS l=0 w=0 x=505716 y=236909 diode_nd2ps_06v0
x a_510063_259404# a_498947_268180# VIN VDD s=816000,16204 d=816000,16204 l=2000 w=8000 x=510063 y=259404 ppolyf_u
x a_499016_248165# VDD s=21168000,22704 l=0 w=0 x=499016 y=248165 diode_pd2nw_06v0
x a_499016_248165# VDD s=21168000,22704 l=0 w=0 x=503448 y=248165 diode_pd2nw_06v0
x a_499016_248165# TEXT$9_0/VSUBS l=0 w=0 x=499020 y=236909 diode_nd2ps_06v0
x a_498947_268180# VDD s=21168000,22704 l=0 w=0 x=498947 y=268180 diode_pd2nw_06v0
x a_498947_268180# TEXT$9_0/VSUBS l=0 w=0 x=498951 y=256924 diode_nd2ps_06v0
x a_499016_248165# VDD s=21168000,22704 l=0 w=0 x=505664 y=248165 diode_pd2nw_06v0
x a_499016_248165# VDD s=21168000,22704 l=0 w=0 x=501232 y=248165 diode_pd2nw_06v0
x a_498947_268180# TEXT$9_0/VSUBS l=0 w=0 x=501183 y=256924 diode_nd2ps_06v0
x a_499016_248165# TEXT$9_0/VSUBS l=0 w=0 x=503484 y=236909 diode_nd2ps_06v0
x a_498947_268180# TEXT$9_0/VSUBS l=0 w=0 x=505647 y=256924 diode_nd2ps_06v0
x a_498947_268180# VDD s=21168000,22704 l=0 w=0 x=503379 y=268180 diode_pd2nw_06v0
x a_510132_239389# a_499016_248165# VBIAS VDD s=816000,16204 d=816000,16204 l=2000 w=8000 x=510132 y=239389 ppolyf_u
x a_499016_248165# TEXT$9_0/VSUBS l=0 w=0 x=501252 y=236909 diode_nd2ps_06v0
x a_498947_268180# TEXT$9_0/VSUBS l=0 w=0 x=503415 y=256924 diode_nd2ps_06v0
C TEXT$23_0/m1_15120_0# TEXT$21_0/m4_15840_0# 0.0
C TEXT$20_0/m3_8640_0# TEXT$3_0/m2_6000_0# 0.0
C TEXT$20_0/m3_6480_0# TEXT$6_0/m4_3600_0# 0.0
C TEXT$20_0/m3_10800_0# TEXT$23_0/m1_10800_0# 0.0
C TEXT$8_0/m4_4800_960# TEXT$9_0/m1_5760_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$3_0/m2_4800_0# 1.1
C TEXT$1_0/m1_12000_0# TEXT$20_0/m3_15120_0# 0.0
C TEXT$6_0/m4_1200_0# TEXT$22_0/m2_3780_0# 0.0
C TEXT$1_0/m1_2400_0# TEXT$4_0/m3_2400_0# 0.0
C M_0/a_403251_244568# VDD 1.1
C TEXT$22_0/m2_8640_0# TEXT$8_0/m4_4800_960# 0.0
C TEXT$1_0/m1_2400_0# TEXT$22_0/m2_4320_0# 0.0
C TEXT$1_0/m1_7200_0# TEXT$6_0/m4_8400_0# 0.0
C TEXT$1_0/m1_8400_0# TEXT$6_0/m4_7200_0# 0.0
C TEXT$7_0/m2_960_0# TEXT$9_0/m1_0_0# 0.0
C TEXT$7_0/m2_0_0# TEXT$9_0/m1_960_0# 0.0
C TEXT$6_0/m4_8400_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$24_0/m3_3840_0# TEXT$23_0/m1_7920_720# 0.0
C TEXT$1_0/m1_9600_0# TEXT$4_0/m3_8400_0# 0.0
C TEXT$4_0/m3_9600_0# TEXT$3_0/m2_9600_0# 1.0
C TEXT$1_0/m1_8400_0# TEXT$4_0/m3_9600_0# 0.0
C TEXT$1_0/m1_8400_0# TEXT$23_0/m1_11700_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$3_0/m2_9600_0# 0.0
C TEXT$23_0/m1_18000_0# TEXT$21_0/m4_18000_0# 0.0
C VDD TEXT$24_0/m3_6720_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$9_0/m1_7680_0# 0.0
C TEXT$20_0/m3_1440_0# TEXT$22_0/m2_720_0# 0.0
C TEXT$23_0/m1_3780_0# TEXT$3_0/m2_1200_0# 0.0
C TEXT$20_0/m3_2160_0# TEXT$22_0/m2_2160_0# 0.4
C TEXT$23_0/m1_15840_0# TEXT$23_0/m1_16560_0# 0.3
C TEXT$6_0/m4_3600_0# TEXT$6_0/m4_4800_0# 0.3
C TEXT$21_0/m4_5760_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$9_0/m1_5760_0# TEXT$7_0/m2_5760_0# 0.7
C TEXT$4_0/m3_6000_0# TEXT$6_0/m4_4800_0# 0.0
C VDD m4_400150_261569# 1.5
C TEXT$21_0/m4_10800_0# TEXT$23_0/m1_10080_0# 0.0
C TEXT$20_0/m3_8640_0# TEXT$9_0/m1_3840_0# 0.0
C TEXT$22_0/m2_9360_0# TEXT$6_0/m4_7200_0# 0.0
C TEXT$4_0/m3_0_0# TEXT$6_0/m4_0_0# 1.1
C M_0/a_402461_244568# VDD 1.2
C TEXT$20_0/m3_720_0# TEXT$23_0/m1_720_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$3_0/m2_2400_0# 0.0
C TEXT$4_0/m3_6000_0# TEXT$4_0/m3_7200_0# 0.3
C TEXT$1_0/m1_6000_0# TEXT$23_0/m1_7920_720# 0.0
C TEXT$7_0/m2_2880_0# TEXT$7_0/m2_3840_0# 0.1
C TEXT$20_0/m3_14400_0# TEXT$3_0/m2_12000_0# 0.0
C TEXT$22_0/m2_17280_0# TEXT$20_0/m3_17280_0# 0.4
C TEXT$8_0/m4_6720_0# TEXT$24_0/m3_6720_0# 0.7
C TEXT$20_0/m3_12960_0# TEXT$22_0/m2_12960_0# 0.4
C TEXT$20_0/m3_17280_0# TEXT$21_0/m4_17280_0# 0.4
C TEXT$1_0/m1_6000_0# TEXT$3_0/m2_6000_0# 1.1
C TEXT$3_0/m2_7200_0# TEXT$3_0/m2_6000_0# 0.3
C TEXT$21_0/m4_10800_0# TEXT$9_0/m1_6720_0# 0.0
C TEXT$24_0/m3_6720_0# TEXT$7_0/m2_6720_0# 0.7
C TEXT$20_0/m3_7200_0# TEXT$8_0/m4_2880_0# 0.0
C TEXT$6_0/m4_1200_0# TEXT$21_0/m4_3780_0# 0.0
C TEXT$24_0/m3_3840_0# TEXT$9_0/m1_3840_0# 0.0
C TEXT$20_0/m3_8640_0# TEXT$8_0/m4_3840_0# 0.0
C TEXT$21_0/m4_7200_0# TEXT$3_0/m2_4800_0# 0.0
C TEXT$1_0/m1_12000_0# TEXT$6_0/m4_12000_0# 0.0
C TEXT$20_0/m3_15120_0# TEXT$20_0/m3_14400_0# 0.3
C TEXT$21_0/m4_9360_0# TEXT$8_0/m4_4800_960# 0.0
C TEXT$20_0/m3_10800_0# TEXT$6_0/m4_8400_0# 0.0
C TEXT$4_0/m3_2400_0# TEXT$22_0/m2_4320_0# 0.0
C m4_400150_261569# m3_419992_265695# 0.1
C VDD M_0/a_395162_259299# 3.1
C TEXT$24_0/m3_7680_0# TEXT$8_0/m4_9600_0# 0.0
C TEXT$4_0/m3_9600_0# TEXT$20_0/m3_11700_0# 0.0
C TEXT$22_0/m2_17280_0# TEXT$22_0/m2_16560_0# 0.1
C TEXT$20_0/m3_3780_0# TEXT$22_0/m2_3780_0# 0.2
C a_498947_268180# VDD 57.0
C TEXT$20_0/m3_720_0# TEXT$21_0/m4_1440_0# 0.0
C TEXT$6_0/m4_4800_0# TEXT$23_0/m1_7200_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$20_0/m3_11700_0# 0.0
C TEXT$22_0/m2_16560_0# TEXT$21_0/m4_17280_0# 0.0
C TEXT$8_0/m4_3840_0# TEXT$24_0/m3_3840_0# 0.7
C TEXT$22_0/m2_11700_0# TEXT$9_0/m1_6720_0# 0.0
C TEXT$20_0/m3_6480_0# TEXT$20_0/m3_7200_0# 0.3
C TEXT$22_0/m2_14400_0# TEXT$8_0/m4_10560_0# 0.0
C TEXT$8_0/m4_2160_0# TEXT$24_0/m3_2880_0# 0.0
C TEXT$20_0/m3_2160_0# TEXT$21_0/m4_2160_0# 0.4
C TEXT$1_0/m1_1200_0# TEXT$3_0/m2_1200_0# 1.1
C TEXT$22_0/m2_10080_0# TEXT$23_0/m1_10800_0# 0.0
C TEXT$8_0/m4_0_0# TEXT$7_0/m2_960_0# 0.0
C TEXT$24_0/m3_0_0# TEXT$7_0/m2_0_0# 0.6
C TEXT$8_0/m4_5760_0# TEXT$7_0/m2_4800_960# 0.0
C TEXT$22_0/m2_5760_0# TEXT$24_0/m3_2160_0# 0.0
C TEXT$24_0/m3_7680_0# TEXT$9_0/m1_6720_0# 0.0
C TEXT$20_0/m3_12960_0# TEXT$21_0/m4_11700_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$21_0/m4_12960_0# 0.0
C TEXT$24_0/m3_960_0# TEXT$7_0/m2_2160_0# 0.0
C TEXT$6_0/m4_7200_0# TEXT$21_0/m4_10080_0# 0.0
C PU EN 0.2
C TEXT$4_0/m3_8400_0# TEXT$21_0/m4_10800_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$22_0/m2_12960_0# 0.0
C VDD M_0/a_383940_262205# 15.5
C M_0/a_395162_259299# m3_419992_265695# 0.0
C TEXT$23_0/m1_4320_0# TEXT$23_0/m1_5760_0# 0.0
C TEXT$20_0/m3_13680_0# TEXT$20_0/m3_14400_0# 0.3
C TEXT$20_0/m3_3780_0# TEXT$22_0/m2_2880_720# 0.0
C TEXT$20_0/m3_2880_720# TEXT$22_0/m2_3780_0# 0.0
C a_498947_268180# m3_419992_265695# 1.7
C M_0/a_404311_244568# VDD 6.4
C TEXT$22_0/m2_7200_0# TEXT$23_0/m1_7920_720# 0.0
C TEXT$20_0/m3_2880_720# TEXT$23_0/m1_2160_0# 0.0
C TEXT$7_0/m2_2160_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$3_0/m2_0_0# TEXT$3_0/m2_1200_0# 0.2
C TEXT$22_0/m2_7920_720# TEXT$3_0/m2_4800_0# 0.0
C TEXT$4_0/m3_6000_0# TEXT$20_0/m3_7920_720# 0.0
C TEXT$20_0/m3_14400_0# TEXT$8_0/m4_9600_0# 0.0
C TEXT$1_0/m1_3600_0# TEXT$4_0/m3_3600_0# 0.0
C VDD TEXT$7_0/m2_960_0# 0.0
C TEXT$1_0/m1_3600_0# TEXT$22_0/m2_5760_0# 0.0
C TEXT$20_0/m3_14400_0# TEXT$6_0/m4_12000_0# 0.0
C TEXT$1_0/m1_9600_0# TEXT$6_0/m4_8400_0# 0.0
C TEXT$21_0/m4_10800_0# TEXT$21_0/m4_11700_0# 0.1
C TEXT$7_0/m2_2160_0# TEXT$9_0/m1_960_0# 0.0
C TEXT$7_0/m2_960_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$6_0/m4_9600_0# TEXT$3_0/m2_9600_0# 0.0
C TEXT$20_0/m3_3780_0# TEXT$21_0/m4_3780_0# 0.2
C TEXT$24_0/m3_7680_0# TEXT$24_0/m3_9600_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$22_0/m2_11700_0# 0.0
C TEXT$1_0/m1_9600_0# TEXT$4_0/m3_10800_0# 0.0
C TEXT$4_0/m3_10800_0# TEXT$3_0/m2_10800_0# 1.2
C TEXT$20_0/m3_15120_0# TEXT$24_0/m3_10560_0# 0.0
C TEXT$22_0/m2_4320_0# TEXT$21_0/m4_5760_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$22_0/m2_10800_0# 0.0
C TEXT$23_0/m1_12960_0# TEXT$3_0/m2_10800_0# 0.0
C TEXT$23_0/m1_8640_0# TEXT$23_0/m1_7920_720# 0.1
C TEXT$21_0/m4_8640_0# TEXT$23_0/m1_7920_720# 0.0
C TEXT$20_0/m3_1440_0# TEXT$22_0/m2_2160_0# 0.0
C M_0/a_383940_262205# m3_419992_265695# 0.0
C TEXT$22_0/m2_0_0# TEXT$22_0/m2_720_0# 0.2
C TEXT$24_0/m3_5760_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$23_0/m1_8640_0# TEXT$3_0/m2_6000_0# 0.0
C TEXT$21_0/m4_10800_0# TEXT$23_0/m1_10800_0# 0.0
C TEXT$21_0/m4_8640_0# TEXT$3_0/m2_6000_0# 0.0
C TEXT$4_0/m3_0_0# TEXT$20_0/m3_2160_0# 0.0
C TEXT$20_0/m3_2880_720# TEXT$22_0/m2_2880_720# 0.2
C M_0/a_404311_244568# m3_419992_265695# 0.3
C M_0/a_403521_244568# VDD 7.5
C TEXT$6_0/m4_4800_0# TEXT$6_0/m4_6000_0# 0.3
C TEXT$21_0/m4_6480_0# TEXT$24_0/m3_2160_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$21_0/m4_11700_0# 0.0
C TEXT$1_0/m1_0_0# TEXT$22_0/m2_2160_0# 0.0
C TEXT$8_0/m4_9600_0# TEXT$9_0/m1_7680_0# 0.0
C TEXT$4_0/m3_7200_0# TEXT$6_0/m4_6000_0# 0.0
C TEXT$20_0/m3_9360_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$4_0/m3_1200_0# TEXT$6_0/m4_1200_0# 1.1
C TEXT$20_0/m3_5760_0# TEXT$3_0/m2_3600_0# 0.0
C TEXT$4_0/m3_7200_0# TEXT$4_0/m3_8400_0# 0.1
C TEXT$22_0/m2_10080_0# TEXT$7_0/m2_5760_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$23_0/m1_7200_0# 0.0
C TEXT$7_0/m2_3840_0# TEXT$7_0/m2_4800_960# 0.1
C TEXT$21_0/m4_11700_0# TEXT$24_0/m3_7680_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$24_0/m3_0_0# 0.0
C TEXT$3_0/m2_1200_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$20_0/m3_3780_0# TEXT$21_0/m4_2880_720# 0.0
C TEXT$20_0/m3_2880_720# TEXT$21_0/m4_3780_0# 0.0
C TEXT$20_0/m3_13680_0# TEXT$22_0/m2_13680_0# 0.3
C TEXT$20_0/m3_18000_0# TEXT$21_0/m4_18000_0# 0.3
C TEXT$8_0/m4_4800_960# TEXT$8_0/m4_5760_0# 0.2
C TEXT$7_0/m2_0_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$23_0/m1_10800_0# 0.0
C TEXT$21_0/m4_7920_720# TEXT$23_0/m1_7920_720# 0.0
C TEXT$9_0/m1_6720_0# TEXT$9_0/m1_7680_0# 0.3
C TEXT$20_0/m3_14400_0# TEXT$24_0/m3_9600_0# 0.0
C TEXT$23_0/m1_3780_0# TEXT$22_0/m2_3780_0# 0.2
C TEXT$6_0/m4_2400_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$24_0/m3_4800_960# TEXT$9_0/m1_4800_960# 0.0
C TEXT$22_0/m2_13680_0# TEXT$8_0/m4_9600_0# 0.0
C TEXT$21_0/m4_7920_720# TEXT$3_0/m2_6000_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$8_0/m4_6720_0# 0.0
C M_0/a_403521_244568# m3_419992_265695# 0.0
C M_0/a_402731_244568# VDD 7.4
C TEXT$1_0/m1_3600_0# TEXT$21_0/m4_6480_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$8_0/m4_2160_0# 0.0
C TEXT$23_0/m1_8640_0# TEXT$9_0/m1_3840_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$6_0/m4_9600_0# 0.0
C TEXT$4_0/m3_3600_0# TEXT$22_0/m2_5760_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$24_0/m3_10560_0# TEXT$8_0/m4_9600_0# 0.0
C TEXT$4_0/m3_10800_0# TEXT$20_0/m3_12960_0# 0.0
C TEXT$6_0/m4_3600_0# TEXT$3_0/m2_3600_0# 0.0
C TEXT$24_0/m3_960_0# TEXT$23_0/m1_5760_0# 0.0
C TEXT$22_0/m2_0_0# TEXT$21_0/m4_720_0# 0.0
C TEXT$20_0/m3_6480_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$20_0/m3_1440_0# TEXT$21_0/m4_2160_0# 0.0
C TEXT$23_0/m1_12960_0# TEXT$20_0/m3_12960_0# 0.0
C TEXT$20_0/m3_7200_0# TEXT$20_0/m3_7920_720# 0.1
C TEXT$20_0/m3_8640_0# TEXT$24_0/m3_3840_0# 0.0
C TEXT$20_0/m3_2880_720# TEXT$21_0/m4_2880_720# 0.2
C TEXT$8_0/m4_5760_0# TEXT$7_0/m2_5760_0# 0.0
C TEXT$22_0/m2_18000_0# TEXT$23_0/m1_18000_0# 0.3
C TEXT$6_0/m4_7200_0# TEXT$23_0/m1_10080_0# 0.0
C TEXT$8_0/m4_960_0# TEXT$7_0/m2_960_0# 0.0
C TEXT$21_0/m4_8640_0# TEXT$8_0/m4_3840_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$24_0/m3_2880_0# 0.0
C TEXT$23_0/m1_15840_0# TEXT$22_0/m2_15840_0# 0.4
C TEXT$24_0/m3_7680_0# TEXT$9_0/m1_9600_0# 0.0
C TEXT$24_0/m3_9600_0# TEXT$9_0/m1_7680_0# 0.0
C TEXT$23_0/m1_4320_0# TEXT$9_0/m1_0_0# 0.0
C TEXT$20_0/m3_13680_0# TEXT$21_0/m4_12960_0# 0.0
C TEXT$20_0/m3_12960_0# TEXT$21_0/m4_13680_0# 0.0
C TEXT$1_0/m1_2400_0# TEXT$6_0/m4_2400_0# 0.0
C TEXT$20_0/m3_15120_0# TEXT$20_0/m3_15840_0# 0.2
C TEXT$23_0/m1_3780_0# TEXT$22_0/m2_2880_720# 0.0
C TEXT$23_0/m1_2880_720# TEXT$22_0/m2_3780_0# 0.0
C VDD M_0/a_374398_259299# 1.8
C TEXT$23_0/m1_6480_0# TEXT$23_0/m1_5760_0# 0.2
C TEXT$20_0/m3_15120_0# TEXT$9_0/m1_10560_0# 0.0
C M_0/a_402731_244568# m3_419992_265695# 0.0
C TEXT$6_0/m4_8400_0# TEXT$21_0/m4_10800_0# 0.0
C M_0/a_401941_244568# VDD 7.4
C TEXT$23_0/m1_2880_720# TEXT$23_0/m1_2160_0# 0.1
C TEXT$23_0/m1_5760_0# TEXT$9_0/m1_960_0# 0.0
C TEXT$22_0/m2_15120_0# TEXT$3_0/m2_12000_0# 0.0
C TEXT$1_0/m1_12000_0# TEXT$22_0/m2_14400_0# 0.0
C TEXT$22_0/m2_12960_0# TEXT$22_0/m2_13680_0# 0.2
C TEXT$4_0/m3_1200_0# TEXT$20_0/m3_3780_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$9_0/m1_6720_0# 0.0
C VDD VIN 19.9
C TEXT$23_0/m1_3780_0# TEXT$21_0/m4_3780_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$6_0/m4_6000_0# 0.0
C TEXT$22_0/m2_13680_0# TEXT$24_0/m3_9600_0# 0.0
C TEXT$1_0/m1_1200_0# TEXT$22_0/m2_3780_0# 0.0
C TEXT$3_0/m2_1200_0# TEXT$3_0/m2_2400_0# 0.3
C TEXT$22_0/m2_10800_0# TEXT$8_0/m4_6720_0# 0.0
C TEXT$9_0/m1_5760_0# TEXT$9_0/m1_4800_960# 0.1
C TEXT$22_0/m2_17280_0# TEXT$21_0/m4_17280_0# 0.0
C TEXT$1_0/m1_4800_0# TEXT$4_0/m3_4800_0# 0.0
C VDD TEXT$7_0/m2_2880_0# 0.0
C TEXT$8_0/m4_4800_960# TEXT$7_0/m2_3840_0# 0.0
C TEXT$20_0/m3_15120_0# TEXT$22_0/m2_15120_0# 0.4
C TEXT$1_0/m1_9600_0# TEXT$6_0/m4_10800_0# 0.0
C TEXT$1_0/m1_10800_0# TEXT$6_0/m4_9600_0# 0.0
C TEXT$7_0/m2_2160_0# TEXT$9_0/m1_2880_0# 0.0
C TEXT$7_0/m2_2880_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$21_0/m4_7920_720# TEXT$8_0/m4_3840_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$6_0/m4_8400_0# 0.0
C TEXT$6_0/m4_10800_0# TEXT$3_0/m2_10800_0# 0.0
C TEXT$22_0/m2_8640_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$22_0/m2_10800_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$21_0/m4_15120_0# TEXT$8_0/m4_10560_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$21_0/m4_4320_0# 0.4
C TEXT$1_0/m1_12000_0# TEXT$4_0/m3_10800_0# 0.0
C TEXT$1_0/m1_10800_0# TEXT$4_0/m3_12000_0# 0.0
C M_0/a_374398_259299# m3_419992_265695# 0.0
C TEXT$24_0/m3_9600_0# TEXT$24_0/m3_10560_0# 0.2
C TEXT$23_0/m1_2880_720# TEXT$22_0/m2_2880_720# 0.2
C TEXT$4_0/m3_3600_0# TEXT$21_0/m4_6480_0# 0.0
C TEXT$4_0/m3_12000_0# TEXT$3_0/m2_12000_0# 1.1
C VDD a_499016_248165# 58.1
C TEXT$21_0/m4_0_0# TEXT$21_0/m4_720_0# 0.2
C TEXT$22_0/m2_5760_0# TEXT$21_0/m4_6480_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$21_0/m4_5760_0# 0.0
C M_0/a_401941_244568# m3_419992_265695# 0.0
C TEXT$23_0/m1_12960_0# TEXT$22_0/m2_11700_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$22_0/m2_12960_0# 0.0
C M_0/a_401151_244568# VDD 44.9
C TEXT$20_0/m3_14400_0# TEXT$9_0/m1_9600_0# 0.0
C TEXT$22_0/m2_720_0# TEXT$22_0/m2_1440_0# 0.2
C TEXT$6_0/m4_6000_0# TEXT$6_0/m4_7200_0# 0.3
C VDD VCM_OUT 0.1
C TEXT$21_0/m4_7200_0# TEXT$24_0/m3_2880_0# 0.0
C TEXT$23_0/m1_2880_720# TEXT$21_0/m4_3780_0# 0.0
C TEXT$4_0/m3_12000_0# TEXT$20_0/m3_15120_0# 0.0
C TEXT$22_0/m2_12960_0# TEXT$21_0/m4_12960_0# 0.0
C TEXT$21_0/m4_14400_0# TEXT$3_0/m2_12000_0# 0.0
C TEXT$4_0/m3_0_0# TEXT$1_0/m1_0_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$6_0/m4_7200_0# 0.0
C TEXT$22_0/m2_4320_0# TEXT$7_0/m2_0_0# 0.0
C TEXT$22_0/m2_720_0# TEXT$23_0/m1_720_0# 0.3
C TEXT$4_0/m3_2400_0# TEXT$6_0/m4_2400_0# 1.0
C TEXT$3_0/m2_0_0# TEXT$23_0/m1_2160_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$4_0/m3_9600_0# 0.3
C TEXT$22_0/m2_4320_0# TEXT$6_0/m4_2400_0# 0.0
C TEXT$1_0/m1_2400_0# TEXT$20_0/m3_4320_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$23_0/m1_11700_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$8_0/m4_960_0# 0.0
C TEXT$20_0/m3_9360_0# TEXT$24_0/m3_5760_0# 0.0
C TEXT$20_0/m3_14400_0# TEXT$22_0/m2_14400_0# 0.4
C a_499016_248165# m3_419992_265695# 0.0
C VDD TEXT$8_0/m4_9600_0# 0.0
C VDD M_0/a_373878_259299# 3.1
C TEXT$20_0/m3_15120_0# TEXT$21_0/m4_14400_0# 0.0
C TEXT$24_0/m3_2160_0# TEXT$7_0/m2_960_0# 0.0
C M_0/a_401151_244568# m3_419992_265695# 2.2
C TEXT$1_0/m1_1200_0# TEXT$21_0/m4_3780_0# 0.0
C TEXT$1_0/m1_6000_0# TEXT$3_0/m2_7200_0# 0.0
C TEXT$9_0/m1_7680_0# TEXT$9_0/m1_9600_0# 0.0
C PU VDD 0.0
C TEXT$4_0/m3_9600_0# TEXT$21_0/m4_11700_0# 0.0
C TEXT$24_0/m3_960_0# TEXT$9_0/m1_0_0# 0.0
C TEXT$8_0/m4_2880_0# TEXT$9_0/m1_2880_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$8_0/m4_7680_0# 0.0
C TEXT$22_0/m2_15120_0# TEXT$6_0/m4_12000_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$21_0/m4_11700_0# 0.0
C VDD BCM_OUT 0.1
C TEXT$23_0/m1_2880_720# TEXT$21_0/m4_2880_720# 0.0
C TEXT$1_0/m1_4800_0# TEXT$21_0/m4_7200_0# 0.0
C VDD TEXT$9_0/m1_6720_0# 0.0
C TEXT$20_0/m3_12960_0# TEXT$6_0/m4_10800_0# 0.0
C TEXT$24_0/m3_4800_960# TEXT$24_0/m3_5760_0# 0.2
C TEXT$21_0/m4_9360_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$22_0/m2_2880_720# TEXT$3_0/m2_0_0# 0.0
C TEXT$6_0/m4_4800_0# TEXT$3_0/m2_4800_0# 0.0
C TEXT$22_0/m2_720_0# TEXT$23_0/m1_1440_0# 0.0
C TEXT$22_0/m2_720_0# TEXT$21_0/m4_1440_0# 0.0
C TEXT$23_0/m1_13680_0# TEXT$20_0/m3_13680_0# 0.0
C TEXT$4_0/m3_6000_0# TEXT$3_0/m2_6000_0# 1.1
C TEXT$21_0/m4_11700_0# TEXT$21_0/m4_12960_0# 0.0
C TEXT$22_0/m2_13680_0# TEXT$9_0/m1_9600_0# 0.0
C M_0/a_403251_244568# M_0/a_404041_244568# 0.3
C TEXT$22_0/m2_3780_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$20_0/m3_9360_0# TEXT$24_0/m3_4800_960# 0.0
C M_0/a_373878_259299# m3_419992_265695# 0.0
C TEXT$23_0/m1_11700_0# TEXT$23_0/m1_10800_0# 0.1
C TEXT$4_0/m3_12000_0# TEXT$6_0/m4_12000_0# 1.1
C TEXT$9_0/m1_0_0# TEXT$9_0/m1_960_0# 0.2
C TEXT$23_0/m1_8640_0# TEXT$20_0/m3_8640_0# 0.0
C TEXT$24_0/m3_9600_0# TEXT$9_0/m1_10560_0# 0.0
C TEXT$24_0/m3_10560_0# TEXT$9_0/m1_9600_0# 0.0
C TEXT$21_0/m4_720_0# TEXT$23_0/m1_720_0# 0.0
C TEXT$20_0/m3_8640_0# TEXT$21_0/m4_8640_0# 0.4
C TEXT$20_0/m3_13680_0# TEXT$21_0/m4_14400_0# 0.0
C TEXT$21_0/m4_720_0# TEXT$23_0/m1_0_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$23_0/m1_3780_0# 0.0
C TEXT$8_0/m4_6720_0# TEXT$9_0/m1_6720_0# 0.0
C TEXT$23_0/m1_16560_0# TEXT$23_0/m1_17280_0# 0.1
C VDD CCM_OUT 0.1
C TEXT$9_0/m1_6720_0# TEXT$7_0/m2_6720_0# 0.7
C TEXT$22_0/m2_13680_0# TEXT$22_0/m2_14400_0# 0.2
C TEXT$8_0/m4_10560_0# TEXT$7_0/m2_10560_0# 0.0
C VDD TEXT$24_0/m3_9600_0# 0.0
C TEXT$21_0/m4_14400_0# TEXT$8_0/m4_9600_0# 0.0
C TEXT$4_0/m3_2400_0# TEXT$20_0/m3_4320_0# 0.0
C TEXT$21_0/m4_14400_0# TEXT$6_0/m4_12000_0# 0.0
C M_0/a_404041_244568# m4_400150_261569# 1.6
C TEXT$21_0/m4_8640_0# TEXT$24_0/m3_3840_0# 0.0
C TEXT$23_0/m1_8640_0# TEXT$24_0/m3_3840_0# 0.0
C TEXT$22_0/m2_4320_0# TEXT$20_0/m3_4320_0# 0.4
C TEXT$22_0/m2_14400_0# TEXT$24_0/m3_10560_0# 0.0
C TEXT$22_0/m2_18000_0# TEXT$20_0/m3_18000_0# 0.3
C M_0/a_402461_244568# M_0/a_404041_244568# 0.1
C TEXT$23_0/m1_7200_0# TEXT$23_0/m1_7920_720# 0.1
C TEXT$20_0/m3_2160_0# TEXT$6_0/m4_0_0# 0.0
C TEXT$3_0/m2_2400_0# TEXT$3_0/m2_3600_0# 0.2
C TEXT$20_0/m3_10080_0# TEXT$3_0/m2_7200_0# 0.0
C VDD TEXT$7_0/m2_4800_960# 0.0
C TEXT$3_0/m2_0_0# TEXT$21_0/m4_2880_720# 0.0
C TEXT$1_0/m1_4800_0# TEXT$22_0/m2_7920_720# 0.0
C TEXT$1_0/m1_12000_0# TEXT$6_0/m4_10800_0# 0.0
C TEXT$7_0/m2_3840_0# TEXT$9_0/m1_2880_0# 0.0
C TEXT$7_0/m2_2880_0# TEXT$9_0/m1_3840_0# 0.0
C TEXT$24_0/m3_5760_0# TEXT$9_0/m1_5760_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$24_0/m3_2160_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$7_0/m2_7680_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$21_0/m4_7200_0# 0.0
C VDD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# 0.2
C TEXT$21_0/m4_720_0# TEXT$21_0/m4_1440_0# 0.3
C TEXT$22_0/m2_6480_0# TEXT$21_0/m4_7200_0# 0.0
C TEXT$1_0/m1_12000_0# TEXT$23_0/m1_14400_0# 0.0
C TEXT$23_0/m1_12960_0# TEXT$22_0/m2_13680_0# 0.0
C TEXT$23_0/m1_13680_0# TEXT$22_0/m2_12960_0# 0.0
C TEXT$23_0/m1_15120_0# TEXT$3_0/m2_12000_0# 0.0
C TEXT$23_0/m1_15840_0# TEXT$21_0/m4_16560_0# 0.0
C TEXT$24_0/m3_7680_0# TEXT$7_0/m2_7680_0# 0.7
C TEXT$22_0/m2_1440_0# TEXT$22_0/m2_2160_0# 0.1
C TEXT$24_0/m3_960_0# TEXT$8_0/m4_0_0# 0.0
C TEXT$8_0/m4_3840_0# TEXT$7_0/m2_2880_0# 0.0
C TEXT$6_0/m4_7200_0# TEXT$6_0/m4_8400_0# 0.1
C TEXT$8_0/m4_2160_0# TEXT$7_0/m2_2160_0# 0.0
C TEXT$23_0/m1_13680_0# TEXT$24_0/m3_9600_0# 0.0
C TEXT$21_0/m4_7920_720# TEXT$24_0/m3_3840_0# 0.0
C TEXT$1_0/m1_6000_0# TEXT$23_0/m1_8640_0# 0.0
C TEXT$20_0/m3_7200_0# TEXT$23_0/m1_7920_720# 0.0
C TEXT$22_0/m2_8640_0# TEXT$20_0/m3_9360_0# 0.0
C TEXT$22_0/m2_13680_0# TEXT$21_0/m4_13680_0# 0.0
C M_0/a_402461_244568# M_0/a_403251_244568# 0.6
C a_498947_268180# M_0/a_404041_244568# 0.6
C TEXT$4_0/m3_8400_0# TEXT$6_0/m4_9600_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$1_0/m1_1200_0# 0.0
C TEXT$4_0/m3_9600_0# TEXT$6_0/m4_8400_0# 0.0
C TEXT$22_0/m2_5760_0# TEXT$7_0/m2_960_0# 0.0
C TEXT$20_0/m3_15120_0# TEXT$23_0/m1_15120_0# 0.0
C TEXT$3_0/m2_3600_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$3_0/m2_4800_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$6_0/m4_8400_0# 0.0
C TEXT$4_0/m3_9600_0# TEXT$4_0/m3_10800_0# 0.2
C TEXT$21_0/m4_14400_0# TEXT$24_0/m3_9600_0# 0.0
C TEXT$21_0/m4_11700_0# TEXT$8_0/m4_6720_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$23_0/m1_12960_0# 0.0
C TEXT$24_0/m3_2880_0# TEXT$7_0/m2_2160_0# 0.0
C TEXT$24_0/m3_2160_0# TEXT$7_0/m2_2880_0# 0.0
C TEXT$20_0/m3_15120_0# TEXT$21_0/m4_15840_0# 0.0
C TEXT$24_0/m3_0_0# TEXT$9_0/m1_0_0# 0.0
C TEXT$22_0/m2_8640_0# TEXT$24_0/m3_4800_960# 0.0
C TEXT$6_0/m4_9600_0# TEXT$21_0/m4_11700_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$21_0/m4_5760_0# 0.0
C VDD VIN_OUT 2.9
C TEXT$9_0/m1_9600_0# TEXT$9_0/m1_10560_0# 0.2
C TEXT$21_0/m4_11700_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$1_0/m1_7200_0# TEXT$3_0/m2_8400_0# 0.0
C VDD TEXT$24_0/m3_960_0# 0.0
C TEXT$4_0/m3_10800_0# TEXT$21_0/m4_12960_0# 0.0
C TEXT$24_0/m3_960_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$6_0/m4_6000_0# TEXT$23_0/m1_7920_720# 0.0
C VDD TEXT$9_0/m1_9600_0# 0.0
C M_0/a_404311_244568# M_0/a_404041_244568# 2.3
C a_498947_268180# M_0/a_403251_244568# 0.6
C TEXT$20_0/m3_13680_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$22_0/m2_7920_720# 0.0
C TEXT$6_0/m4_6000_0# TEXT$3_0/m2_6000_0# 0.0
C TEXT$22_0/m2_2160_0# TEXT$23_0/m1_1440_0# 0.0
C TEXT$8_0/m4_9600_0# TEXT$8_0/m4_7680_0# 0.0
C TEXT$23_0/m1_10800_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$22_0/m2_1440_0# TEXT$21_0/m4_2160_0# 0.0
C TEXT$21_0/m4_9360_0# TEXT$24_0/m3_5760_0# 0.0
C TEXT$23_0/m1_14400_0# TEXT$20_0/m3_14400_0# 0.0
C TEXT$21_0/m4_12960_0# TEXT$21_0/m4_13680_0# 0.2
C TEXT$22_0/m2_14400_0# TEXT$9_0/m1_10560_0# 0.0
C TEXT$1_0/m1_3600_0# TEXT$6_0/m4_3600_0# 0.0
C VDD M_0/a_365708_259299# 48.9
C TEXT$8_0/m4_4800_960# VDD 0.0
C TEXT$23_0/m1_6480_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$20_0/m3_3780_0# TEXT$6_0/m4_1200_0# 0.0
C VDD TEXT$9_0/m1_960_0# 0.0
C TEXT$8_0/m4_9600_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$8_0/m4_2880_0# TEXT$8_0/m4_2160_0# 0.2
C TEXT$3_0/m2_1200_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$22_0/m2_9360_0# TEXT$3_0/m2_7200_0# 0.0
C TEXT$9_0/m1_960_0# TEXT$9_0/m1_2160_0# 0.1
C TEXT$20_0/m3_9360_0# TEXT$21_0/m4_9360_0# 0.4
C TEXT$20_0/m3_14400_0# TEXT$21_0/m4_15120_0# 0.0
C TEXT$23_0/m1_15120_0# TEXT$6_0/m4_12000_0# 0.0
C M_0/a_395162_259299# m4_400150_261569# 0.9
C a_498947_268180# m4_400150_261569# 0.1
C TEXT$23_0/m1_17280_0# TEXT$23_0/m1_18000_0# 0.2
C TEXT$9_0/m1_7680_0# TEXT$7_0/m2_7680_0# 0.7
C M_0/a_404311_244568# M_0/a_403251_244568# 0.1
C a_498947_268180# M_0/a_402461_244568# 0.6
C M_0/a_403521_244568# M_0/a_404041_244568# 2.4
C TEXT$22_0/m2_14400_0# TEXT$22_0/m2_15120_0# 0.2
C TEXT$8_0/m4_2880_0# TEXT$24_0/m3_2880_0# 0.7
C TEXT$20_0/m3_6480_0# TEXT$8_0/m4_2160_0# 0.0
C TEXT$22_0/m2_2160_0# TEXT$23_0/m1_2160_0# 0.4
C TEXT$4_0/m3_3600_0# TEXT$20_0/m3_5760_0# 0.0
C TEXT$23_0/m1_13680_0# TEXT$9_0/m1_9600_0# 0.0
C TEXT$21_0/m4_9360_0# TEXT$24_0/m3_4800_960# 0.0
C TEXT$22_0/m2_5760_0# TEXT$20_0/m3_5760_0# 0.4
C M_0/a_365708_259299# m3_419992_265695# 0.7
C VDD TEXT$7_0/m2_5760_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$3_0/m2_3600_0# TEXT$3_0/m2_4800_0# 0.3
C TEXT$20_0/m3_10800_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$23_0/m1_8640_0# TEXT$21_0/m4_8640_0# 0.0
C TEXT$1_0/m1_0_0# TEXT$6_0/m4_0_0# 0.0
C TEXT$7_0/m2_3840_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$20_0/m3_6480_0# TEXT$24_0/m3_2880_0# 0.0
C TEXT$21_0/m4_2160_0# TEXT$23_0/m1_1440_0# 0.0
C TEXT$4_0/m3_12000_0# TEXT$22_0/m2_14400_0# 0.0
C TEXT$8_0/m4_0_0# TEXT$24_0/m3_0_0# 0.6
C TEXT$24_0/m3_9600_0# TEXT$8_0/m4_7680_0# 0.0
C TEXT$23_0/m1_17280_0# TEXT$20_0/m3_16560_0# 0.0
C TEXT$23_0/m1_16560_0# TEXT$20_0/m3_17280_0# 0.0
C TEXT$22_0/m2_4320_0# TEXT$23_0/m1_5760_0# 0.0
C M_0/a_383940_262205# m4_400150_261569# 0.5
C TEXT$21_0/m4_1440_0# TEXT$21_0/m4_2160_0# 0.1
C TEXT$22_0/m2_7200_0# TEXT$21_0/m4_7920_720# 0.0
C TEXT$22_0/m2_10080_0# TEXT$24_0/m3_5760_0# 0.0
C TEXT$23_0/m1_14400_0# TEXT$22_0/m2_13680_0# 0.0
C M_0/a_402731_244568# M_0/a_404041_244568# 0.2
C M_0/a_404311_244568# M_0/a_402461_244568# 0.1
C M_0/a_403521_244568# M_0/a_403251_244568# 2.3
C TEXT$22_0/m2_2160_0# TEXT$22_0/m2_2880_720# 0.1
C TEXT$24_0/m3_9600_0# TEXT$7_0/m2_9600_0# 0.7
C TEXT$24_0/m3_960_0# TEXT$8_0/m4_960_0# 0.7
C TEXT$8_0/m4_6720_0# TEXT$7_0/m2_5760_0# 0.0
C TEXT$4_0/m3_3600_0# TEXT$6_0/m4_3600_0# 1.1
C TEXT$4_0/m3_6000_0# TEXT$20_0/m3_8640_0# 0.0
C TEXT$22_0/m2_5760_0# TEXT$6_0/m4_3600_0# 0.0
C TEXT$6_0/m4_8400_0# TEXT$6_0/m4_9600_0# 0.3
C TEXT$23_0/m1_14400_0# TEXT$24_0/m3_10560_0# 0.0
C TEXT$21_0/m4_10080_0# TEXT$3_0/m2_7200_0# 0.0
C TEXT$22_0/m2_10080_0# TEXT$20_0/m3_9360_0# 0.0
C TEXT$22_0/m2_9360_0# TEXT$20_0/m3_10080_0# 0.0
C TEXT$22_0/m2_14400_0# TEXT$21_0/m4_14400_0# 0.0
C TEXT$4_0/m3_9600_0# TEXT$6_0/m4_10800_0# 0.0
C TEXT$4_0/m3_10800_0# TEXT$6_0/m4_9600_0# 0.0
C TEXT$7_0/m2_5760_0# TEXT$7_0/m2_6720_0# 0.2
C TEXT$22_0/m2_6480_0# TEXT$7_0/m2_2160_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$22_0/m2_8640_0# 0.1
C TEXT$4_0/m3_10800_0# TEXT$4_0/m3_12000_0# 0.1
C TEXT$21_0/m4_7920_720# TEXT$21_0/m4_8640_0# 0.1
C TEXT$23_0/m1_11700_0# TEXT$7_0/m2_7680_0# 0.0
C TEXT$23_0/m1_16560_0# TEXT$22_0/m2_16560_0# 0.4
C TEXT$21_0/m4_15120_0# TEXT$24_0/m3_10560_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$24_0/m3_6720_0# 0.0
C TEXT$21_0/m4_11700_0# TEXT$8_0/m4_7680_0# 0.0
C TEXT$20_0/m3_15840_0# TEXT$20_0/m3_16560_0# 0.3
C VDD TEXT$24_0/m3_0_0# 0.0
C M_0/a_383940_262205# M_0/a_395162_259299# 1.0
C TEXT$23_0/m1_12960_0# TEXT$23_0/m1_13680_0# 0.2
C TEXT$24_0/m3_3840_0# TEXT$7_0/m2_2880_0# 0.0
C TEXT$8_0/m4_960_0# TEXT$9_0/m1_960_0# 0.0
C TEXT$6_0/m4_10800_0# TEXT$21_0/m4_12960_0# 0.0
C TEXT$20_0/m3_6480_0# TEXT$21_0/m4_5760_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$21_0/m4_6480_0# 0.0
C TEXT$1_0/m1_9600_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$1_0/m1_8400_0# TEXT$3_0/m2_9600_0# 0.0
C M_0/a_403521_244568# M_0/a_402461_244568# 0.1
C M_0/a_402731_244568# M_0/a_403251_244568# 2.4
C M_0/a_401941_244568# M_0/a_404041_244568# 0.2
C M_0/a_404311_244568# a_498947_268180# 0.6
C TEXT$8_0/m4_5760_0# TEXT$24_0/m3_5760_0# 0.7
C TEXT$22_0/m2_8640_0# TEXT$21_0/m4_9360_0# 0.0
C TEXT$23_0/m1_13680_0# TEXT$21_0/m4_13680_0# 0.0
C TEXT$20_0/m3_14400_0# TEXT$7_0/m2_10560_0# 0.0
C TEXT$20_0/m3_2880_720# TEXT$20_0/m3_3780_0# 0.1
C TEXT$22_0/m2_4320_0# TEXT$3_0/m2_1200_0# 0.0
C TEXT$22_0/m2_18000_0# TEXT$21_0/m4_18000_0# 0.0
C PU PD 0.4
C TEXT$20_0/m3_4320_0# TEXT$7_0/m2_0_0# 0.0
C TEXT$20_0/m3_15840_0# TEXT$22_0/m2_15840_0# 0.4
C TEXT$22_0/m2_2160_0# TEXT$21_0/m4_2880_720# 0.0
C TEXT$21_0/m4_13680_0# TEXT$21_0/m4_14400_0# 0.3
C TEXT$1_0/m1_4800_0# TEXT$6_0/m4_4800_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$6_0/m4_2400_0# 0.0
C VDD TEXT$9_0/m1_2880_0# 0.0
C TEXT$8_0/m4_4800_960# TEXT$9_0/m1_3840_0# 0.0
C TEXT$1_0/m1_6000_0# TEXT$4_0/m3_6000_0# 0.0
C M_0/a_403251_244568# M_0/a_410724_251737# 1.5
C TEXT$1_0/m1_7200_0# TEXT$22_0/m2_10080_0# 0.0
C TEXT$6_0/m4_3600_0# TEXT$21_0/m4_6480_0# 0.0
C TEXT$9_0/m1_2160_0# TEXT$9_0/m1_2880_0# 0.1
C TEXT$20_0/m3_10080_0# TEXT$21_0/m4_10080_0# 0.4
C M_0/a_403521_244568# a_498947_268180# 0.6
C M_0/a_401151_244568# M_0/a_404041_244568# 0.6
C M_0/a_401941_244568# M_0/a_403251_244568# 0.2
C M_0/a_402731_244568# M_0/a_402461_244568# 2.3
C TEXT$8_0/m4_7680_0# TEXT$9_0/m1_9600_0# 0.0
C TEXT$8_0/m4_0_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$3_0/m2_7200_0# TEXT$23_0/m1_9360_0# 0.0
C TEXT$20_0/m3_1440_0# TEXT$20_0/m3_2160_0# 0.1
C TEXT$22_0/m2_15120_0# TEXT$22_0/m2_15840_0# 0.2
C TEXT$9_0/m1_9600_0# TEXT$7_0/m2_9600_0# 0.7
C TEXT$22_0/m2_10800_0# TEXT$24_0/m3_6720_0# 0.0
C TEXT$24_0/m3_960_0# TEXT$24_0/m3_2160_0# 0.1
C TEXT$8_0/m4_4800_960# TEXT$8_0/m4_3840_0# 0.2
C TEXT$4_0/m3_0_0# TEXT$23_0/m1_2160_0# 0.0
C TEXT$23_0/m1_14400_0# TEXT$9_0/m1_10560_0# 0.0
C TEXT$3_0/m2_4800_0# TEXT$23_0/m1_7920_720# 0.0
C TEXT$22_0/m2_10080_0# TEXT$9_0/m1_5760_0# 0.0
C TEXT$1_0/m1_0_0# TEXT$20_0/m3_2160_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$20_0/m3_6480_0# 0.4
C TEXT$22_0/m2_4320_0# TEXT$9_0/m1_0_0# 0.0
C VDD TEXT$7_0/m2_7680_0# 0.0
C TEXT$1_0/m1_8400_0# TEXT$20_0/m3_11700_0# 0.0
C TEXT$3_0/m2_4800_0# TEXT$3_0/m2_6000_0# 0.2
C TEXT$20_0/m3_10080_0# TEXT$22_0/m2_10800_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$3_0/m2_9600_0# 0.0
C TEXT$22_0/m2_5760_0# TEXT$23_0/m1_4320_0# 0.0
C M_0/a_403251_244568# M_0/a_410134_251737# 1.9
C M_0/a_383620_262205# M_0/a_383940_262205# 1.1
C TEXT$24_0/m3_2160_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$22_0/m2_3780_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$1_0/m1_1200_0# TEXT$6_0/m4_1200_0# 0.0
C TEXT$1_0/m1_2400_0# TEXT$3_0/m2_3600_0# 0.0
C TEXT$21_0/m4_15120_0# TEXT$9_0/m1_10560_0# 0.0
C TEXT$22_0/m2_14400_0# TEXT$7_0/m2_9600_0# 0.0
C M_0/a_403521_244568# M_0/a_404311_244568# 0.8
C M_0/a_401151_244568# M_0/a_403251_244568# 0.1
C M_0/a_401941_244568# M_0/a_402461_244568# 2.4
C M_0/a_402731_244568# a_498947_268180# 0.6
C TEXT$24_0/m3_2160_0# TEXT$9_0/m1_960_0# 0.0
C TEXT$8_0/m4_960_0# TEXT$24_0/m3_0_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$23_0/m1_5760_0# 0.0
C TEXT$23_0/m1_18000_0# TEXT$20_0/m3_17280_0# 0.0
C TEXT$21_0/m4_2160_0# TEXT$21_0/m4_2880_720# 0.2
C TEXT$23_0/m1_14400_0# TEXT$22_0/m2_15120_0# 0.0
C TEXT$3_0/m2_7200_0# TEXT$23_0/m1_10080_0# 0.0
C TEXT$23_0/m1_15120_0# TEXT$22_0/m2_14400_0# 0.0
C TEXT$23_0/m1_3780_0# TEXT$20_0/m3_3780_0# 0.0
C TEXT$4_0/m3_0_0# TEXT$22_0/m2_2880_720# 0.0
C TEXT$24_0/m3_10560_0# TEXT$7_0/m2_10560_0# 0.7
C TEXT$20_0/m3_8640_0# TEXT$6_0/m4_6000_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$6_0/m4_4800_0# 1.1
C TEXT$4_0/m3_7200_0# TEXT$20_0/m3_9360_0# 0.0
C sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# PD 0.0
C TEXT$6_0/m4_9600_0# TEXT$6_0/m4_10800_0# 0.2
C TEXT$20_0/m3_8640_0# TEXT$7_0/m2_4800_960# 0.0
C TEXT$21_0/m4_10800_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$21_0/m4_7200_0# TEXT$8_0/m4_2880_0# 0.0
C TEXT$22_0/m2_10080_0# TEXT$20_0/m3_10800_0# 0.0
C TEXT$22_0/m2_15120_0# TEXT$21_0/m4_15120_0# 0.0
C TEXT$4_0/m3_12000_0# TEXT$6_0/m4_10800_0# 0.0
C TEXT$7_0/m2_6720_0# TEXT$7_0/m2_7680_0# 0.2
C TEXT$22_0/m2_7200_0# TEXT$7_0/m2_2880_0# 0.0
C TEXT$8_0/m4_5760_0# TEXT$9_0/m1_5760_0# 0.0
C M_0/a_404041_244568# M_0/a_409498_256643# 0.9
C TEXT$6_0/m4_0_0# TEXT$3_0/m2_1200_0# 0.0
C TEXT$1_0/m1_3600_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$1_0/m1_4800_0# TEXT$20_0/m3_7920_720# 0.0
C M_0/a_401941_244568# a_498947_268180# 2.9
C M_0/a_401151_244568# M_0/a_402461_244568# 0.1
C M_0/a_402731_244568# M_0/a_404311_244568# 0.3
C TEXT$20_0/m3_16560_0# TEXT$20_0/m3_17280_0# 0.1
C TEXT$23_0/m1_13680_0# TEXT$23_0/m1_14400_0# 0.3
C TEXT$24_0/m3_4800_960# TEXT$7_0/m2_3840_0# 0.0
C TEXT$24_0/m3_3840_0# TEXT$7_0/m2_4800_960# 0.0
C TEXT$23_0/m1_2880_720# TEXT$20_0/m3_3780_0# 0.0
C TEXT$23_0/m1_3780_0# TEXT$20_0/m3_2880_720# 0.0
C TEXT$20_0/m3_6480_0# TEXT$21_0/m4_7200_0# 0.0
C TEXT$1_0/m1_8400_0# TEXT$22_0/m2_10800_0# 0.0
C TEXT$1_0/m1_9600_0# TEXT$3_0/m2_10800_0# 0.0
C TEXT$1_0/m1_10800_0# TEXT$3_0/m2_9600_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$4_0/m3_12000_0# TEXT$21_0/m4_15120_0# 0.0
C TEXT$4_0/m3_6000_0# TEXT$23_0/m1_8640_0# 0.0
C TEXT$4_0/m3_6000_0# TEXT$21_0/m4_8640_0# 0.0
C M_0/a_403251_244568# BCM_OUT 0.2
C M_0/a_404041_244568# CCM_OUT 0.0
C M_0/a_402461_244568# VCM_OUT 0.2
C TEXT$21_0/m4_3780_0# TEXT$21_0/m4_4320_0# 0.1
C TEXT$22_0/m2_10080_0# TEXT$21_0/m4_9360_0# 0.0
C TEXT$22_0/m2_9360_0# TEXT$21_0/m4_10080_0# 0.0
C M_0/a_377450_262205# M_0/a_383620_262205# 0.5
C M_0/a_374398_259299# M_0/a_383940_262205# 0.3
C TEXT$23_0/m1_8640_0# TEXT$23_0/m1_9360_0# 0.3
C TEXT$20_0/m3_5760_0# TEXT$7_0/m2_960_0# 0.0
C TEXT$20_0/m3_16560_0# TEXT$22_0/m2_16560_0# 0.4
C TEXT$4_0/m3_0_0# TEXT$21_0/m4_2880_720# 0.0
C TEXT$22_0/m2_7200_0# TEXT$23_0/m1_7200_0# 0.4
C a_498947_268180# a_499016_248165# 0.1
C TEXT$21_0/m4_14400_0# TEXT$21_0/m4_15120_0# 0.3
C TEXT$24_0/m3_6720_0# TEXT$9_0/m1_6720_0# 0.0
C TEXT$20_0/m3_10080_0# TEXT$23_0/m1_10080_0# 0.0
C TEXT$1_0/m1_6000_0# TEXT$6_0/m4_6000_0# 0.0
C TEXT$6_0/m4_6000_0# TEXT$3_0/m2_7200_0# 0.0
C TEXT$22_0/m2_4320_0# TEXT$8_0/m4_0_0# 0.0
C M_0/a_401941_244568# M_0/a_404311_244568# 0.3
C M_0/a_402731_244568# M_0/a_403521_244568# 0.8
C M_0/a_401151_244568# a_498947_268180# 3.4
C VDD TEXT$9_0/m1_4800_960# 0.0
C TEXT$22_0/m2_17280_0# TEXT$23_0/m1_16560_0# 0.0
C TEXT$4_0/m3_7200_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$1_0/m1_7200_0# TEXT$4_0/m3_7200_0# 0.0
C TEXT$9_0/m1_2880_0# TEXT$9_0/m1_3840_0# 0.1
C TEXT$22_0/m2_5760_0# TEXT$24_0/m3_960_0# 0.0
C TEXT$6_0/m4_1200_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$23_0/m1_2880_720# TEXT$20_0/m3_2880_720# 0.0
C TEXT$6_0/m4_4800_0# TEXT$21_0/m4_7200_0# 0.0
C TEXT$23_0/m1_16560_0# TEXT$21_0/m4_17280_0# 0.0
C TEXT$20_0/m3_10800_0# TEXT$21_0/m4_10800_0# 0.4
C TEXT$20_0/m3_0_0# TEXT$22_0/m2_0_0# 0.4
C TEXT$4_0/m3_6000_0# TEXT$21_0/m4_7920_720# 0.0
C TEXT$22_0/m2_15840_0# TEXT$22_0/m2_16560_0# 0.2
C TEXT$9_0/m1_10560_0# TEXT$7_0/m2_10560_0# 0.7
C TEXT$4_0/m3_3600_0# TEXT$23_0/m1_6480_0# 0.0
C m4_400150_261569# M_0/a_409498_256643# 3.3
C VDD TEXT$8_0/m4_2160_0# 0.0
C TEXT$20_0/m3_8640_0# TEXT$8_0/m4_4800_960# 0.0
C TEXT$22_0/m2_4320_0# TEXT$22_0/m2_3780_0# 0.1
C TEXT$22_0/m2_5760_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$20_0/m3_7920_720# 0.0
C M_0/a_404041_244568# M_0/a_409618_260539# 3.0
C M_0/a_374398_259299# M_0/a_383620_262205# 0.9
C TEXT$8_0/m4_2160_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$22_0/m2_7200_0# TEXT$20_0/m3_7200_0# 0.4
C TEXT$22_0/m2_8640_0# TEXT$7_0/m2_3840_0# 0.0
C VDD TEXT$7_0/m2_10560_0# 0.0
C M_0/a_401941_244568# M_0/a_403521_244568# 0.3
C M_0/a_401151_244568# M_0/a_404311_244568# 2.4
C TEXT$20_0/m3_10800_0# TEXT$22_0/m2_11700_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$22_0/m2_10800_0# 0.0
C TEXT$20_0/m3_12960_0# TEXT$3_0/m2_10800_0# 0.0
C TEXT$20_0/m3_15840_0# TEXT$21_0/m4_16560_0# 0.0
C TEXT$1_0/m1_3600_0# TEXT$3_0/m2_4800_0# 0.0
C TEXT$22_0/m2_15120_0# TEXT$7_0/m2_10560_0# 0.0
C m4_400150_261569# CCM_OUT 0.6
C VDD TEXT$24_0/m3_2880_0# 0.0
C TEXT$8_0/m4_4800_960# TEXT$24_0/m3_3840_0# 0.0
C TEXT$24_0/m3_2160_0# TEXT$9_0/m1_2880_0# 0.0
C TEXT$24_0/m3_2880_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$22_0/m2_9360_0# TEXT$23_0/m1_9360_0# 0.4
C M_0/a_404041_244568# VIN_OUT 2.5
C TEXT$21_0/m4_5760_0# TEXT$3_0/m2_3600_0# 0.0
C VDD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# 0.3
C TEXT$21_0/m4_7920_720# TEXT$23_0/m1_7200_0# 0.0
C TEXT$4_0/m3_0_0# TEXT$4_0/m3_1200_0# 0.3
C TEXT$20_0/m3_9360_0# TEXT$6_0/m4_7200_0# 0.0
C TEXT$8_0/m4_7680_0# TEXT$7_0/m2_7680_0# 0.0
C M_0/a_374398_259299# M_0/a_377450_262205# 36.6
C TEXT$20_0/m3_2880_720# TEXT$3_0/m2_0_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$6_0/m4_4800_0# 0.0
C TEXT$22_0/m2_10800_0# TEXT$21_0/m4_10080_0# 0.0
C TEXT$21_0/m4_11700_0# TEXT$24_0/m3_6720_0# 0.0
C TEXT$20_0/m3_0_0# TEXT$21_0/m4_0_0# 0.4
C TEXT$22_0/m2_15840_0# TEXT$21_0/m4_15840_0# 0.0
C TEXT$7_0/m2_7680_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$7_0/m2_3840_0# 0.0
C M_0/a_401941_244568# M_0/a_402731_244568# 0.8
C M_0/a_401151_244568# M_0/a_403521_244568# 1.5
C TEXT$23_0/m1_2880_720# TEXT$23_0/m1_3780_0# 0.1
C TEXT$4_0/m3_1200_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$6_0/m4_1200_0# TEXT$3_0/m2_2400_0# 0.0
C TEXT$23_0/m1_14400_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$20_0/m3_3780_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$22_0/m2_10080_0# TEXT$8_0/m4_5760_0# 0.0
C TEXT$20_0/m3_17280_0# TEXT$20_0/m3_18000_0# 0.2
C TEXT$22_0/m2_9360_0# TEXT$23_0/m1_10080_0# 0.0
C M_0/a_403251_244568# VIN_OUT 0.1
C TEXT$23_0/m1_14400_0# TEXT$23_0/m1_15120_0# 0.3
C TEXT$8_0/m4_2880_0# TEXT$7_0/m2_2160_0# 0.0
C TEXT$21_0/m4_6480_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$23_0/m1_5760_0# 0.0
C TEXT$24_0/m3_6720_0# TEXT$23_0/m1_10800_0# 0.0
C TEXT$6_0/m4_6000_0# TEXT$21_0/m4_8640_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$21_0/m4_7200_0# 0.0
C TEXT$20_0/m3_7200_0# TEXT$21_0/m4_7920_720# 0.0
C TEXT$21_0/m4_14400_0# TEXT$7_0/m2_10560_0# 0.0
C TEXT$1_0/m1_9600_0# TEXT$22_0/m2_11700_0# 0.0
C TEXT$1_0/m1_12000_0# TEXT$3_0/m2_10800_0# 0.0
C TEXT$1_0/m1_10800_0# TEXT$3_0/m2_12000_0# 0.0
C TEXT$4_0/m3_7200_0# TEXT$21_0/m4_9360_0# 0.0
C m4_400150_261569# M_0/a_409618_260539# 3.6
C TEXT$21_0/m4_8640_0# TEXT$7_0/m2_4800_960# 0.0
C TEXT$23_0/m1_8640_0# TEXT$7_0/m2_4800_960# 0.0
C TEXT$22_0/m2_10080_0# TEXT$21_0/m4_10800_0# 0.0
C TEXT$1_0/m1_1200_0# TEXT$23_0/m1_3780_0# 0.0
C TEXT$23_0/m1_15120_0# TEXT$21_0/m4_15120_0# 0.0
C TEXT$20_0/m3_10080_0# TEXT$23_0/m1_10800_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$6_0/m4_3600_0# 0.0
C M_0/a_401151_244568# M_0/a_402731_244568# 1.5
C TEXT$22_0/m2_6480_0# TEXT$3_0/m2_3600_0# 0.0
C TEXT$20_0/m3_6480_0# TEXT$7_0/m2_2160_0# 0.0
C TEXT$8_0/m4_2160_0# TEXT$8_0/m4_960_0# 0.2
C TEXT$20_0/m3_15120_0# TEXT$3_0/m2_12000_0# 0.0
C TEXT$1_0/m1_7200_0# TEXT$6_0/m4_7200_0# 0.0
C TEXT$21_0/m4_15120_0# TEXT$21_0/m4_15840_0# 0.2
C TEXT$7_0/m2_0_0# TEXT$9_0/m1_0_0# 0.6
C TEXT$6_0/m4_7200_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$6_0/m4_0_0# TEXT$23_0/m1_2160_0# 0.0
C m4_400150_261569# VIN_OUT 0.2
C TEXT$4_0/m3_9600_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$22_0/m2_17280_0# TEXT$23_0/m1_18000_0# 0.0
C TEXT$1_0/m1_8400_0# TEXT$4_0/m3_8400_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$3_0/m2_9600_0# 0.0
C M_0/a_402461_244568# VIN_OUT 0.1
C TEXT$9_0/m1_3840_0# TEXT$9_0/m1_4800_960# 0.1
C TEXT$23_0/m1_11700_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$23_0/m1_17280_0# TEXT$21_0/m4_18000_0# 0.0
C TEXT$6_0/m4_6000_0# TEXT$21_0/m4_7920_720# 0.0
C M_0/a_410134_251737# M_0/a_410724_251737# 0.4
C VDD TEXT$24_0/m3_5760_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$9_0/m1_6720_0# 0.0
C TEXT$20_0/m3_720_0# TEXT$22_0/m2_720_0# 0.3
C TEXT$20_0/m3_14400_0# TEXT$8_0/m4_10560_0# 0.0
C a_499016_248165# M_0/a_374398_259299# 0.5
C TEXT$20_0/m3_2160_0# TEXT$22_0/m2_1440_0# 0.0
C TEXT$21_0/m4_11700_0# TEXT$3_0/m2_9600_0# 0.0
C TEXT$1_0/m1_8400_0# TEXT$21_0/m4_11700_0# 0.0
C M_0/a_401151_244568# M_0/a_401941_244568# 1.8
C TEXT$6_0/m4_0_0# TEXT$22_0/m2_2880_720# 0.0
C TEXT$20_0/m3_0_0# TEXT$23_0/m1_0_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$3_0/m2_1200_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$20_0/m3_7920_720# 0.2
C TEXT$1_0/m1_4800_0# TEXT$23_0/m1_7920_720# 0.0
C TEXT$4_0/m3_7200_0# TEXT$22_0/m2_10080_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$22_0/m2_9360_0# TEXT$7_0/m2_4800_960# 0.0
C TEXT$22_0/m2_17280_0# TEXT$20_0/m3_16560_0# 0.0
C TEXT$20_0/m3_12960_0# TEXT$22_0/m2_11700_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$22_0/m2_12960_0# 0.0
C TEXT$20_0/m3_17280_0# TEXT$21_0/m4_16560_0# 0.0
C TEXT$20_0/m3_16560_0# TEXT$21_0/m4_17280_0# 0.0
C a_498947_268180# VIN_OUT 0.5
C TEXT$1_0/m1_4800_0# TEXT$3_0/m2_6000_0# 0.0
C TEXT$1_0/m1_8400_0# TEXT$23_0/m1_10800_0# 0.0
C VDD TEXT$24_0/m3_4800_960# 0.0
C TEXT$24_0/m3_6720_0# TEXT$7_0/m2_5760_0# 0.0
C TEXT$1_0/m1_2400_0# TEXT$1_0/m1_3600_0# 0.2
C TEXT$24_0/m3_3840_0# TEXT$9_0/m1_2880_0# 0.0
C TEXT$23_0/m1_2880_720# TEXT$3_0/m2_0_0# 0.0
C TEXT$3_0/m2_12000_0# TEXT$6_0/m4_12000_0# 0.0
C M_0/a_373878_259299# M_0/a_374398_259299# 0.9
C TEXT$22_0/m2_10800_0# TEXT$23_0/m1_10080_0# 0.0
C TEXT$21_0/m4_8640_0# TEXT$8_0/m4_4800_960# 0.0
C TEXT$4_0/m3_1200_0# TEXT$4_0/m3_2400_0# 0.3
C TEXT$21_0/m4_5760_0# TEXT$8_0/m4_960_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$22_0/m2_4320_0# 0.0
C TEXT$20_0/m3_10080_0# TEXT$7_0/m2_5760_0# 0.0
C TEXT$23_0/m1_3780_0# TEXT$23_0/m1_4320_0# 0.1
C TEXT$4_0/m3_8400_0# TEXT$20_0/m3_11700_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$21_0/m4_10800_0# 0.0
C M_0/a_410724_251737# BCM_OUT 1.2
C TEXT$23_0/m1_11700_0# TEXT$20_0/m3_10800_0# 0.0
C TEXT$20_0/m3_720_0# TEXT$21_0/m4_720_0# 0.3
C TEXT$22_0/m2_16560_0# TEXT$21_0/m4_16560_0# 0.0
C TEXT$22_0/m2_10800_0# TEXT$9_0/m1_6720_0# 0.0
C TEXT$7_0/m2_9600_0# TEXT$7_0/m2_10560_0# 0.1
C TEXT$20_0/m3_15120_0# TEXT$6_0/m4_12000_0# 0.0
C TEXT$8_0/m4_2160_0# TEXT$24_0/m3_2160_0# 0.4
C TEXT$20_0/m3_2160_0# TEXT$21_0/m4_1440_0# 0.0
C TEXT$1_0/m1_0_0# TEXT$3_0/m2_1200_0# 0.0
C M_0/a_404311_244568# VIN_OUT 2.4
C TEXT$20_0/m3_4320_0# TEXT$9_0/m1_0_0# 0.0
C TEXT$7_0/m2_2880_0# TEXT$23_0/m1_7200_0# 0.0
C TEXT$6_0/m4_2400_0# TEXT$3_0/m2_3600_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$23_0/m1_15120_0# TEXT$7_0/m2_10560_0# 0.0
C TEXT$8_0/m4_0_0# TEXT$7_0/m2_0_0# 0.0
C TEXT$22_0/m2_5760_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$21_0/m4_11700_0# 0.2
C TEXT$24_0/m3_10560_0# TEXT$8_0/m4_10560_0# 0.8
C TEXT$6_0/m4_0_0# TEXT$21_0/m4_2880_720# 0.0
C VDD M_0/a_386992_259299# 48.8
C TEXT$24_0/m3_960_0# TEXT$7_0/m2_960_0# 0.7
C TEXT$8_0/m4_2880_0# TEXT$7_0/m2_3840_0# 0.0
C M_0/a_373878_259299# a_499016_248165# 1.0
C TEXT$6_0/m4_7200_0# TEXT$21_0/m4_9360_0# 0.0
C TEXT$1_0/m1_10800_0# TEXT$22_0/m2_12960_0# 0.0
C TEXT$24_0/m3_2160_0# TEXT$24_0/m3_2880_0# 0.1
C TEXT$23_0/m1_10080_0# TEXT$23_0/m1_9360_0# 0.1
C TEXT$4_0/m3_4800_0# TEXT$23_0/m1_7920_720# 0.0
C M_0/a_410134_251737# BCM_OUT 0.1
C TEXT$20_0/m3_11700_0# TEXT$23_0/m1_10800_0# 0.0
C VDD TEXT$9_0/m1_5760_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$24_0/m3_7680_0# 0.0
C TEXT$20_0/m3_2160_0# TEXT$23_0/m1_2160_0# 0.0
C TEXT$22_0/m2_7200_0# TEXT$3_0/m2_4800_0# 0.0
C M_0/a_403521_244568# VIN_OUT 0.1
C TEXT$20_0/m3_13680_0# TEXT$8_0/m4_9600_0# 0.0
C TEXT$20_0/m3_7200_0# TEXT$7_0/m2_2880_0# 0.0
C TEXT$1_0/m1_2400_0# TEXT$4_0/m3_3600_0# 0.0
C VDD TEXT$7_0/m2_0_0# 0.0
C TEXT$22_0/m2_9360_0# TEXT$8_0/m4_4800_960# 0.0
C TEXT$1_0/m1_8400_0# TEXT$6_0/m4_8400_0# 0.0
C TEXT$21_0/m4_15840_0# TEXT$21_0/m4_16560_0# 0.3
C TEXT$7_0/m2_960_0# TEXT$9_0/m1_960_0# 0.7
C TEXT$6_0/m4_9600_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$6_0/m4_8400_0# TEXT$3_0/m2_9600_0# 0.0
C TEXT$1_0/m1_1200_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$22_0/m2_10800_0# 0.0
C TEXT$1_0/m1_9600_0# TEXT$4_0/m3_9600_0# 0.0
C TEXT$4_0/m3_10800_0# TEXT$3_0/m2_9600_0# 0.0
C TEXT$4_0/m3_9600_0# TEXT$3_0/m2_10800_0# 0.0
C M_0/a_386992_259299# m3_419992_265695# 0.8
C TEXT$1_0/m1_9600_0# TEXT$23_0/m1_11700_0# 0.0
C TEXT$20_0/m3_1440_0# TEXT$22_0/m2_1440_0# 0.4
C TEXT$20_0/m3_2880_720# TEXT$22_0/m2_2160_0# 0.0
C TEXT$21_0/m4_5760_0# TEXT$24_0/m3_2160_0# 0.0
C TEXT$22_0/m2_10800_0# TEXT$21_0/m4_11700_0# 0.0
C TEXT$21_0/m4_12960_0# TEXT$3_0/m2_10800_0# 0.0
C TEXT$4_0/m3_6000_0# TEXT$6_0/m4_6000_0# 1.1
C M_0/a_402731_244568# VIN_OUT 0.1
C TEXT$20_0/m3_8640_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$22_0/m2_10080_0# TEXT$6_0/m4_7200_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$6_0/m4_0_0# 0.0
C TEXT$20_0/m3_7200_0# TEXT$23_0/m1_7200_0# 0.0
C TEXT$22_0/m2_7200_0# TEXT$9_0/m1_2880_0# 0.0
C TEXT$22_0/m2_17280_0# TEXT$20_0/m3_18000_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$8_0/m4_0_0# 0.0
C TEXT$20_0/m3_12960_0# TEXT$22_0/m2_13680_0# 0.0
C TEXT$20_0/m3_13680_0# TEXT$22_0/m2_12960_0# 0.0
C TEXT$20_0/m3_18000_0# TEXT$21_0/m4_17280_0# 0.0
C TEXT$20_0/m3_17280_0# TEXT$21_0/m4_18000_0# 0.0
C TEXT$22_0/m2_10800_0# TEXT$23_0/m1_10800_0# 0.4
C TEXT$20_0/m3_5760_0# TEXT$24_0/m3_960_0# 0.0
C TEXT$7_0/m2_4800_960# TEXT$23_0/m1_9360_0# 0.0
C TEXT$1_0/m1_3600_0# TEXT$1_0/m1_4800_0# 0.3
C TEXT$8_0/m4_10560_0# TEXT$9_0/m1_10560_0# 0.0
C TEXT$20_0/m3_13680_0# TEXT$24_0/m3_9600_0# 0.0
C TEXT$6_0/m4_1200_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$24_0/m3_4800_960# TEXT$9_0/m1_3840_0# 0.0
C TEXT$24_0/m3_3840_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$21_0/m4_7920_720# TEXT$3_0/m2_4800_0# 0.0
C TEXT$20_0/m3_10800_0# TEXT$8_0/m4_6720_0# 0.0
C TEXT$23_0/m1_15840_0# TEXT$20_0/m3_15840_0# 0.0
C TEXT$4_0/m3_2400_0# TEXT$4_0/m3_3600_0# 0.2
C TEXT$20_0/m3_11700_0# TEXT$6_0/m4_8400_0# 0.0
C TEXT$20_0/m3_10800_0# TEXT$7_0/m2_6720_0# 0.0
C VDD TEXT$8_0/m4_10560_0# 0.0
C TEXT$24_0/m3_9600_0# TEXT$8_0/m4_9600_0# 0.7
C TEXT$20_0/m3_4320_0# TEXT$22_0/m2_3780_0# 0.0
C M_0/a_401941_244568# VIN_OUT 0.1
C TEXT$22_0/m2_4320_0# TEXT$22_0/m2_5760_0# 0.0
C TEXT$20_0/m3_1440_0# TEXT$23_0/m1_1440_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$22_0/m2_0_0# TEXT$21_0/m4_0_0# 0.0
C sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# PD 0.0
C TEXT$23_0/m1_11700_0# TEXT$20_0/m3_12960_0# 0.0
C TEXT$20_0/m3_1440_0# TEXT$21_0/m4_1440_0# 0.4
C TEXT$23_0/m1_12960_0# TEXT$20_0/m3_11700_0# 0.0
C TEXT$8_0/m4_3840_0# TEXT$24_0/m3_4800_960# 0.0
C TEXT$22_0/m2_11700_0# TEXT$9_0/m1_7680_0# 0.0
C TEXT$22_0/m2_15120_0# TEXT$8_0/m4_10560_0# 0.0
C TEXT$20_0/m3_2160_0# TEXT$21_0/m4_2880_720# 0.0
C TEXT$20_0/m3_2880_720# TEXT$21_0/m4_2160_0# 0.0
C TEXT$1_0/m1_1200_0# TEXT$3_0/m2_2400_0# 0.0
C TEXT$22_0/m2_8640_0# TEXT$3_0/m2_6000_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$9_0/m1_960_0# 0.0
C TEXT$22_0/m2_18000_0# TEXT$23_0/m1_17280_0# 0.0
C TEXT$8_0/m4_960_0# TEXT$7_0/m2_0_0# 0.0
C TEXT$24_0/m3_0_0# TEXT$7_0/m2_960_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$24_0/m3_2160_0# 0.0
C TEXT$23_0/m1_15840_0# TEXT$22_0/m2_15120_0# 0.0
C TEXT$24_0/m3_7680_0# TEXT$9_0/m1_7680_0# 0.0
C TEXT$20_0/m3_12960_0# TEXT$21_0/m4_12960_0# 0.4
C TEXT$1_0/m1_2400_0# TEXT$6_0/m4_1200_0# 0.0
C M_0/a_365708_259299# M_0/a_374398_259299# 0.1
C TEXT$21_0/m4_10080_0# TEXT$7_0/m2_5760_0# 0.0
C M_0/a_409498_256643# CCM_OUT 2.2
C TEXT$22_0/m2_14400_0# TEXT$3_0/m2_12000_0# 0.0
C TEXT$24_0/m3_2880_0# TEXT$24_0/m3_3840_0# 0.1
C M_0/a_401151_244568# VIN_OUT 1.0
C PU sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# 0.0
C TEXT$20_0/m3_1440_0# TEXT$23_0/m1_2160_0# 0.0
C TEXT$6_0/m4_3600_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$23_0/m1_7920_720# 0.2
C TEXT$20_0/m3_7920_720# TEXT$6_0/m4_4800_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$3_0/m2_6000_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$7_0/m2_3840_0# 0.0
C TEXT$22_0/m2_17280_0# TEXT$21_0/m4_16560_0# 0.0
C TEXT$1_0/m1_3600_0# TEXT$4_0/m3_4800_0# 0.0
C VDD TEXT$7_0/m2_2160_0# 0.0
C TEXT$1_0/m1_0_0# TEXT$23_0/m1_2160_0# 0.0
C TEXT$20_0/m3_15120_0# TEXT$22_0/m2_14400_0# 0.0
C TEXT$1_0/m1_3600_0# TEXT$22_0/m2_6480_0# 0.0
C TEXT$1_0/m1_9600_0# TEXT$6_0/m4_9600_0# 0.0
C TEXT$21_0/m4_16560_0# TEXT$21_0/m4_17280_0# 0.2
C TEXT$7_0/m2_2160_0# TEXT$9_0/m1_2160_0# 0.3
C TEXT$22_0/m2_10800_0# TEXT$6_0/m4_8400_0# 0.0
C TEXT$6_0/m4_10800_0# TEXT$3_0/m2_9600_0# 0.0
C TEXT$6_0/m4_9600_0# TEXT$3_0/m2_10800_0# 0.0
C TEXT$22_0/m2_8640_0# TEXT$9_0/m1_3840_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$21_0/m4_3780_0# 0.0
C TEXT$21_0/m4_6480_0# TEXT$8_0/m4_2160_0# 0.0
C TEXT$21_0/m4_14400_0# TEXT$8_0/m4_10560_0# 0.0
C TEXT$20_0/m3_3780_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$1_0/m1_10800_0# TEXT$4_0/m3_10800_0# 0.0
C M_0/a_365708_259299# a_499016_248165# 29.5
C TEXT$23_0/m1_2880_720# TEXT$22_0/m2_2160_0# 0.0
C TEXT$4_0/m3_3600_0# TEXT$21_0/m4_5760_0# 0.0
C TEXT$4_0/m3_9600_0# TEXT$22_0/m2_11700_0# 0.0
C TEXT$4_0/m3_12000_0# TEXT$3_0/m2_10800_0# 0.0
C TEXT$23_0/m1_10800_0# TEXT$23_0/m1_10080_0# 0.3
C TEXT$22_0/m2_5760_0# TEXT$21_0/m4_5760_0# 0.0
C TEXT$1_0/m1_10800_0# TEXT$23_0/m1_12960_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$22_0/m2_11700_0# 0.2
C TEXT$20_0/m3_13680_0# TEXT$9_0/m1_9600_0# 0.0
C TEXT$4_0/m3_0_0# TEXT$20_0/m3_2880_720# 0.0
C TEXT$22_0/m2_8640_0# TEXT$8_0/m4_3840_0# 0.0
C TEXT$23_0/m1_10800_0# TEXT$9_0/m1_6720_0# 0.0
C TEXT$21_0/m4_6480_0# TEXT$24_0/m3_2880_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$24_0/m3_7680_0# 0.0
C TEXT$22_0/m2_12960_0# TEXT$21_0/m4_11700_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$21_0/m4_12960_0# 0.0
C M_0/a_409618_260539# M_0/a_409498_256643# 0.4
C TEXT$1_0/m1_0_0# TEXT$22_0/m2_2880_720# 0.0
C TEXT$4_0/m3_7200_0# TEXT$6_0/m4_7200_0# 0.7
C TEXT$8_0/m4_9600_0# TEXT$9_0/m1_9600_0# 0.0
C TEXT$22_0/m2_0_0# TEXT$23_0/m1_0_0# 0.4
C TEXT$22_0/m2_0_0# TEXT$23_0/m1_720_0# 0.0
C TEXT$20_0/m3_6480_0# TEXT$3_0/m2_3600_0# 0.0
C TEXT$4_0/m3_2400_0# TEXT$6_0/m4_1200_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$6_0/m4_2400_0# 0.0
C TEXT$23_0/m1_6480_0# TEXT$23_0/m1_7200_0# 0.3
C TEXT$22_0/m2_4320_0# TEXT$6_0/m4_1200_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$9_0/m1_3840_0# 0.0
C TEXT$3_0/m2_2400_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$20_0/m3_14400_0# TEXT$22_0/m2_13680_0# 0.0
C M_0/a_365708_259299# M_0/a_373878_259299# 1.0
C VDD TEXT$8_0/m4_5760_0# 0.0
C M_0/a_409618_260539# CCM_OUT 0.0
C TEXT$1_0/m1_4800_0# TEXT$1_0/m1_6000_0# 0.2
C TEXT$8_0/m4_2880_0# VDD 0.0
C TEXT$20_0/m3_14400_0# TEXT$24_0/m3_10560_0# 0.0
C TEXT$3_0/m2_3600_0# TEXT$23_0/m1_5760_0# 0.0
C TEXT$22_0/m2_14400_0# TEXT$8_0/m4_9600_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$21_0/m4_11700_0# 0.0
C TEXT$20_0/m3_8640_0# TEXT$20_0/m3_9360_0# 0.3
C TEXT$22_0/m2_14400_0# TEXT$6_0/m4_12000_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$8_0/m4_3840_0# 0.0
C TEXT$4_0/m3_3600_0# TEXT$4_0/m3_4800_0# 0.3
C TEXT$23_0/m1_8640_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$21_0/m4_8640_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$22_0/m2_2160_0# TEXT$3_0/m2_0_0# 0.0
C TEXT$4_0/m3_3600_0# TEXT$22_0/m2_6480_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$7_0/m2_7680_0# 0.0
C TEXT$6_0/m4_3600_0# TEXT$3_0/m2_4800_0# 0.0
C TEXT$22_0/m2_5760_0# TEXT$22_0/m2_6480_0# 0.2
C TEXT$8_0/m4_5760_0# TEXT$8_0/m4_6720_0# 0.2
C TEXT$22_0/m2_720_0# TEXT$21_0/m4_720_0# 0.0
C TEXT$21_0/m4_5760_0# TEXT$21_0/m4_6480_0# 0.2
C TEXT$23_0/m1_13680_0# TEXT$20_0/m3_12960_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$23_0/m1_10800_0# 0.0
C TEXT$20_0/m3_8640_0# TEXT$24_0/m3_4800_960# 0.0
C TEXT$20_0/m3_6480_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$23_0/m1_10080_0# TEXT$7_0/m2_5760_0# 0.0
C TEXT$22_0/m2_7200_0# TEXT$24_0/m3_2880_0# 0.0
C TEXT$4_0/m3_10800_0# TEXT$6_0/m4_12000_0# 0.0
C TEXT$24_0/m3_9600_0# TEXT$9_0/m1_9600_0# 0.0
C TEXT$21_0/m4_10800_0# TEXT$8_0/m4_6720_0# 0.0
C TEXT$20_0/m3_13680_0# TEXT$21_0/m4_13680_0# 0.3
C TEXT$1_0/m1_3600_0# TEXT$6_0/m4_2400_0# 0.0
C TEXT$21_0/m4_11700_0# TEXT$23_0/m1_10800_0# 0.0
C TEXT$21_0/m4_10800_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$1_0/m1_12000_0# TEXT$22_0/m2_15120_0# 0.0
C TEXT$9_0/m1_6720_0# TEXT$7_0/m2_5760_0# 0.0
C TEXT$24_0/m3_3840_0# TEXT$24_0/m3_4800_960# 0.2
C VDD TEXT$24_0/m3_7680_0# 0.0
C TEXT$8_0/m4_10560_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$21_0/m4_13680_0# TEXT$8_0/m4_9600_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$20_0/m3_4320_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$9_0/m1_7680_0# 0.0
C TEXT$22_0/m2_4320_0# TEXT$20_0/m3_3780_0# 0.0
C VDD VBIAS 19.6
C TEXT$23_0/m1_15120_0# TEXT$8_0/m4_10560_0# 0.0
C TEXT$23_0/m1_3780_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$22_0/m2_14400_0# TEXT$24_0/m3_9600_0# 0.0
C TEXT$22_0/m2_18000_0# TEXT$20_0/m3_17280_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$8_0/m4_6720_0# 0.0
C TEXT$20_0/m3_9360_0# TEXT$3_0/m2_7200_0# 0.0
C TEXT$22_0/m2_17280_0# TEXT$21_0/m4_18000_0# 0.0
C TEXT$8_0/m4_4800_960# TEXT$7_0/m2_4800_960# 0.0
C VDD TEXT$7_0/m2_3840_0# 0.0
C TEXT$3_0/m2_4800_0# TEXT$23_0/m1_7200_0# 0.0
C TEXT$23_0/m1_15840_0# TEXT$23_0/m1_15120_0# 0.2
C TEXT$1_0/m1_4800_0# TEXT$22_0/m2_7200_0# 0.0
C TEXT$1_0/m1_10800_0# TEXT$6_0/m4_10800_0# 0.0
C TEXT$21_0/m4_17280_0# TEXT$21_0/m4_18000_0# 0.2
C TEXT$7_0/m2_2880_0# TEXT$9_0/m1_2880_0# 0.7
C TEXT$3_0/m2_0_0# TEXT$21_0/m4_2160_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$6_0/m4_9600_0# 0.0
C TEXT$6_0/m4_10800_0# TEXT$3_0/m2_12000_0# 0.0
C M_0/a_409618_260539# VIN_OUT 0.0
C TEXT$22_0/m2_9360_0# TEXT$9_0/m1_4800_960# 0.0
C VDD EN 20.7
C TEXT$22_0/m2_11700_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$1_0/m1_12000_0# TEXT$4_0/m3_12000_0# 0.0
C TEXT$6_0/m4_0_0# TEXT$6_0/m4_1200_0# 0.3
C TEXT$4_0/m3_10800_0# TEXT$22_0/m2_12960_0# 0.0
C TEXT$24_0/m3_7680_0# TEXT$8_0/m4_6720_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$21_0/m4_6480_0# 0.0
C TEXT$23_0/m1_12960_0# TEXT$22_0/m2_12960_0# 0.4
C TEXT$23_0/m1_14400_0# TEXT$3_0/m2_12000_0# 0.0
C TEXT$23_0/m1_15840_0# TEXT$21_0/m4_15840_0# 0.0
C TEXT$24_0/m3_7680_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$20_0/m3_14400_0# TEXT$9_0/m1_10560_0# 0.0
C TEXT$8_0/m4_2160_0# TEXT$7_0/m2_960_0# 0.0
C TEXT$22_0/m2_13680_0# TEXT$21_0/m4_12960_0# 0.0
C TEXT$22_0/m2_8640_0# TEXT$20_0/m3_8640_0# 0.4
C TEXT$22_0/m2_12960_0# TEXT$21_0/m4_13680_0# 0.0
C TEXT$21_0/m4_15120_0# TEXT$3_0/m2_12000_0# 0.0
C TEXT$24_0/m3_5760_0# TEXT$24_0/m3_6720_0# 0.2
C TEXT$22_0/m2_3780_0# TEXT$3_0/m2_1200_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$1_0/m1_0_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$6_0/m4_8400_0# 1.1
C TEXT$20_0/m3_7200_0# TEXT$3_0/m2_4800_0# 0.0
C TEXT$4_0/m3_3600_0# TEXT$6_0/m4_2400_0# 0.0
C TEXT$7_0/m2_4800_960# TEXT$7_0/m2_5760_0# 0.1
C TEXT$21_0/m4_13680_0# TEXT$24_0/m3_9600_0# 0.0
C TEXT$20_0/m3_10080_0# TEXT$24_0/m3_5760_0# 0.0
C TEXT$20_0/m3_14400_0# TEXT$22_0/m2_15120_0# 0.0
C TEXT$23_0/m1_7200_0# TEXT$9_0/m1_2880_0# 0.0
C TEXT$24_0/m3_2160_0# TEXT$7_0/m2_2160_0# 0.3
C TEXT$20_0/m3_15120_0# TEXT$21_0/m4_15120_0# 0.4
C TEXT$8_0/m4_0_0# TEXT$9_0/m1_0_0# 0.0
C TEXT$22_0/m2_8640_0# TEXT$24_0/m3_3840_0# 0.0
C TEXT$1_0/m1_1200_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$6_0/m4_8400_0# TEXT$21_0/m4_11700_0# 0.0
C TEXT$24_0/m3_0_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$1_0/m1_7200_0# TEXT$3_0/m2_7200_0# 0.7
C TEXT$1_0/m1_6000_0# TEXT$1_0/m1_7200_0# 0.3
C TEXT$23_0/m1_0_0# TEXT$23_0/m1_720_0# 0.3
C TEXT$3_0/m2_7200_0# TEXT$3_0/m2_8400_0# 0.1
C TEXT$24_0/m3_960_0# TEXT$9_0/m1_960_0# 0.0
C TEXT$8_0/m4_2880_0# TEXT$9_0/m1_3840_0# 0.0
C TEXT$20_0/m3_9360_0# TEXT$20_0/m3_10080_0# 0.1
C TEXT$23_0/m1_11700_0# TEXT$21_0/m4_12960_0# 0.0
C TEXT$1_0/m1_4800_0# TEXT$21_0/m4_7920_720# 0.0
C TEXT$6_0/m4_4800_0# TEXT$23_0/m1_7920_720# 0.0
C VDD TEXT$9_0/m1_7680_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$20_0/m3_8640_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$22_0/m2_7200_0# 0.0
C TEXT$4_0/m3_0_0# TEXT$3_0/m2_0_0# 1.1
C TEXT$7_0/m2_3840_0# TEXT$23_0/m1_7920_720# 0.0
C TEXT$4_0/m3_12000_0# TEXT$20_0/m3_14400_0# 0.0
C TEXT$6_0/m4_4800_0# TEXT$3_0/m2_6000_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$22_0/m2_7200_0# 0.2
C TEXT$22_0/m2_1440_0# TEXT$23_0/m1_1440_0# 0.4
C TEXT$22_0/m2_1440_0# TEXT$21_0/m4_1440_0# 0.0
C TEXT$21_0/m4_6480_0# TEXT$21_0/m4_7200_0# 0.3
C TEXT$22_0/m2_14400_0# TEXT$9_0/m1_9600_0# 0.0
C TEXT$8_0/m4_2880_0# TEXT$8_0/m4_3840_0# 0.2
C VDD TEXT$9_0/m1_0_0# 0.0
C TEXT$20_0/m3_7200_0# TEXT$9_0/m1_2880_0# 0.0
C TEXT$8_0/m4_9600_0# TEXT$7_0/m2_7680_0# 0.0
C TEXT$6_0/m4_10800_0# TEXT$6_0/m4_12000_0# 0.1
C TEXT$22_0/m2_7920_720# TEXT$24_0/m3_3840_0# 0.0
C TEXT$1_0/m1_6000_0# TEXT$22_0/m2_8640_0# 0.0
C TEXT$1_0/m1_2400_0# TEXT$1_0/m1_1200_0# 0.3
C TEXT$3_0/m2_1200_0# TEXT$21_0/m4_3780_0# 0.0
C TEXT$23_0/m1_1440_0# TEXT$23_0/m1_720_0# 0.3
C TEXT$24_0/m3_10560_0# TEXT$9_0/m1_10560_0# 0.0
C TEXT$21_0/m4_1440_0# TEXT$23_0/m1_720_0# 0.0
C TEXT$20_0/m3_8640_0# TEXT$21_0/m4_9360_0# 0.0
C TEXT$20_0/m3_14400_0# TEXT$21_0/m4_14400_0# 0.4
C TEXT$21_0/m4_5760_0# TEXT$7_0/m2_960_0# 0.0
C TEXT$22_0/m2_4320_0# TEXT$23_0/m1_3780_0# 0.0
C TEXT$9_0/m1_7680_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$8_0/m4_2880_0# TEXT$24_0/m3_2160_0# 0.0
C VDD TEXT$24_0/m3_10560_0# 0.0
C TEXT$22_0/m2_1440_0# TEXT$23_0/m1_2160_0# 0.0
C TEXT$21_0/m4_15120_0# TEXT$6_0/m4_12000_0# 0.0
C TEXT$22_0/m2_5760_0# TEXT$20_0/m3_4320_0# 0.0
C TEXT$21_0/m4_8640_0# TEXT$24_0/m3_4800_960# 0.0
C TEXT$23_0/m1_8640_0# TEXT$24_0/m3_4800_960# 0.0
C TEXT$22_0/m2_4320_0# TEXT$20_0/m3_5760_0# 0.0
C TEXT$22_0/m2_15120_0# TEXT$24_0/m3_10560_0# 0.0
C TEXT$8_0/m4_4800_960# TEXT$7_0/m2_5760_0# 0.0
C TEXT$20_0/m3_2880_720# TEXT$6_0/m4_0_0# 0.0
C TEXT$1_0/m1_7200_0# TEXT$20_0/m3_10080_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$8_0/m4_7680_0# 0.0
C M_0/a_386992_259299# m4_400150_261569# 0.1
C TEXT$1_0/m1_6000_0# TEXT$22_0/m2_7920_720# 0.0
C TEXT$7_0/m2_3840_0# TEXT$9_0/m1_3840_0# 0.7
C TEXT$21_0/m4_13680_0# TEXT$9_0/m1_9600_0# 0.0
C TEXT$22_0/m2_12960_0# TEXT$6_0/m4_10800_0# 0.0
C TEXT$24_0/m3_6720_0# TEXT$9_0/m1_5760_0# 0.0
C TEXT$20_0/m3_6480_0# TEXT$24_0/m3_2160_0# 0.0
C TEXT$6_0/m4_1200_0# TEXT$6_0/m4_2400_0# 0.3
C TEXT$21_0/m4_1440_0# TEXT$23_0/m1_1440_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$21_0/m4_7920_720# 0.0
C TEXT$24_0/m3_7680_0# TEXT$8_0/m4_7680_0# 0.7
C TEXT$23_0/m1_16560_0# TEXT$20_0/m3_16560_0# 0.0
C TEXT$22_0/m2_7200_0# TEXT$21_0/m4_7200_0# 0.0
C TEXT$1_0/m1_12000_0# TEXT$23_0/m1_15120_0# 0.0
C TEXT$22_0/m2_9360_0# TEXT$24_0/m3_5760_0# 0.0
C TEXT$23_0/m1_13680_0# TEXT$22_0/m2_13680_0# 0.3
C TEXT$23_0/m1_9360_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$24_0/m3_7680_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$24_0/m3_9600_0# TEXT$7_0/m2_7680_0# 0.0
C TEXT$20_0/m3_10080_0# TEXT$9_0/m1_5760_0# 0.0
C TEXT$24_0/m3_960_0# TEXT$24_0/m3_0_0# 0.2
C TEXT$8_0/m4_3840_0# TEXT$7_0/m2_3840_0# 0.0
C TEXT$24_0/m3_2160_0# TEXT$23_0/m1_5760_0# 0.0
C TEXT$20_0/m3_15120_0# TEXT$7_0/m2_10560_0# 0.0
C TEXT$8_0/m4_2160_0# TEXT$7_0/m2_2880_0# 0.0
C TEXT$23_0/m1_14400_0# TEXT$24_0/m3_9600_0# 0.0
C TEXT$21_0/m4_9360_0# TEXT$3_0/m2_7200_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$23_0/m1_7920_720# 0.0
C TEXT$22_0/m2_9360_0# TEXT$20_0/m3_9360_0# 0.4
C TEXT$22_0/m2_13680_0# TEXT$21_0/m4_14400_0# 0.0
C TEXT$4_0/m3_2400_0# TEXT$1_0/m1_1200_0# 0.0
C TEXT$4_0/m3_9600_0# TEXT$6_0/m4_9600_0# 1.0
C TEXT$1_0/m1_1200_0# TEXT$22_0/m2_4320_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$3_0/m2_6000_0# 0.0
C M_0/a_386992_259299# M_0/a_395162_259299# 1.0
C TEXT$23_0/m1_11700_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$23_0/m1_16560_0# TEXT$22_0/m2_15840_0# 0.0
C TEXT$23_0/m1_2160_0# TEXT$23_0/m1_1440_0# 0.1
C TEXT$21_0/m4_14400_0# TEXT$24_0/m3_10560_0# 0.0
C TEXT$1_0/m1_3600_0# TEXT$20_0/m3_6480_0# 0.0
C TEXT$20_0/m3_10800_0# TEXT$24_0/m3_6720_0# 0.0
C VDD TEXT$8_0/m4_0_0# 0.0
C TEXT$24_0/m3_2880_0# TEXT$7_0/m2_2880_0# 0.7
C TEXT$24_0/m3_0_0# TEXT$9_0/m1_960_0# 0.0
C TEXT$22_0/m2_9360_0# TEXT$24_0/m3_4800_960# 0.0
C TEXT$1_0/m1_2400_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$21_0/m4_5760_0# 0.4
C TEXT$1_0/m1_8400_0# TEXT$3_0/m2_8400_0# 1.1
C TEXT$1_0/m1_7200_0# TEXT$1_0/m1_8400_0# 0.1
C TEXT$3_0/m2_8400_0# TEXT$3_0/m2_9600_0# 0.2
C TEXT$22_0/m2_8640_0# TEXT$21_0/m4_8640_0# 0.0
C TEXT$22_0/m2_8640_0# TEXT$23_0/m1_8640_0# 0.4
C TEXT$20_0/m3_10080_0# TEXT$20_0/m3_10800_0# 0.2
C TEXT$1_0/m1_3600_0# TEXT$23_0/m1_5760_0# 0.0
C TEXT$23_0/m1_12960_0# TEXT$21_0/m4_13680_0# 0.0
C VDD TEXT$9_0/m1_10560_0# 0.0
C TEXT$22_0/m2_17280_0# TEXT$22_0/m2_18000_0# 0.2
C TEXT$20_0/m3_14400_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$3_0/m2_1200_0# 1.1
C TEXT$22_0/m2_18000_0# TEXT$21_0/m4_17280_0# 0.0
C M_0/a_386992_259299# M_0/a_383940_262205# 29.5
C TEXT$22_0/m2_7200_0# TEXT$22_0/m2_7920_720# 0.1
C TEXT$20_0/m3_15840_0# TEXT$22_0/m2_15120_0# 0.0
C TEXT$22_0/m2_2160_0# TEXT$21_0/m4_2160_0# 0.0
C TEXT$21_0/m4_7200_0# TEXT$21_0/m4_7920_720# 0.1
C TEXT$21_0/m4_10080_0# TEXT$24_0/m3_5760_0# 0.0
C TEXT$23_0/m1_15120_0# TEXT$20_0/m3_14400_0# 0.0
C TEXT$22_0/m2_15120_0# TEXT$9_0/m1_10560_0# 0.0
C TEXT$1_0/m1_4800_0# TEXT$6_0/m4_3600_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$6_0/m4_1200_0# 0.0
C VDD TEXT$9_0/m1_2160_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$9_0/m1_3840_0# 0.0
C TEXT$8_0/m4_9600_0# TEXT$7_0/m2_10560_0# 0.0
C TEXT$1_0/m1_4800_0# TEXT$4_0/m3_6000_0# 0.0
C TEXT$1_0/m1_7200_0# TEXT$22_0/m2_9360_0# 0.0
C TEXT$3_0/m2_2400_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$6_0/m4_3600_0# TEXT$21_0/m4_5760_0# 0.0
C TEXT$22_0/m2_10080_0# TEXT$3_0/m2_7200_0# 0.0
C TEXT$24_0/m3_2880_0# TEXT$23_0/m1_7200_0# 0.0
C TEXT$20_0/m3_9360_0# TEXT$21_0/m4_10080_0# 0.0
C TEXT$8_0/m4_7680_0# TEXT$9_0/m1_7680_0# 0.0
C TEXT$21_0/m4_6480_0# TEXT$7_0/m2_2160_0# 0.0
C TEXT$20_0/m3_0_0# TEXT$20_0/m3_720_0# 0.2
C TEXT$22_0/m2_7920_720# TEXT$23_0/m1_8640_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$21_0/m4_8640_0# 0.0
C TEXT$23_0/m1_2880_720# TEXT$6_0/m4_0_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$8_0/m4_3840_0# 0.0
C TEXT$9_0/m1_7680_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$9_0/m1_9600_0# TEXT$7_0/m2_7680_0# 0.0
C TEXT$22_0/m2_2880_720# TEXT$22_0/m2_3780_0# 0.1
C TEXT$8_0/m4_2880_0# TEXT$24_0/m3_3840_0# 0.0
C TEXT$20_0/m3_2160_0# TEXT$20_0/m3_2880_720# 0.1
C VDD TEXT$8_0/m4_6720_0# 0.0
C TEXT$4_0/m3_3600_0# TEXT$20_0/m3_6480_0# 0.0
C TEXT$23_0/m1_14400_0# TEXT$9_0/m1_9600_0# 0.0
C PU sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# 0.0
C TEXT$22_0/m2_5760_0# TEXT$20_0/m3_6480_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$20_0/m3_5760_0# 0.0
C VDD m3_419992_265695# 60.5
C TEXT$7_0/m2_0_0# TEXT$7_0/m2_960_0# 0.2
C VDD TEXT$7_0/m2_6720_0# 0.0
C TEXT$4_0/m3_2400_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$22_0/m2_4320_0# TEXT$23_0/m1_4320_0# 0.4
C TEXT$22_0/m2_8640_0# TEXT$22_0/m2_9360_0# 0.2
C TEXT$23_0/m1_8640_0# TEXT$21_0/m4_9360_0# 0.0
C TEXT$21_0/m4_8640_0# TEXT$21_0/m4_9360_0# 0.3
C TEXT$22_0/m2_3780_0# TEXT$21_0/m4_3780_0# 0.0
C TEXT$1_0/m1_1200_0# TEXT$6_0/m4_0_0# 0.0
C TEXT$1_0/m1_2400_0# TEXT$3_0/m2_2400_0# 1.0
C TEXT$7_0/m2_4800_960# TEXT$9_0/m1_4800_960# 0.4
C TEXT$21_0/m4_14400_0# TEXT$9_0/m1_10560_0# 0.0
C TEXT$20_0/m3_7200_0# TEXT$24_0/m3_2880_0# 0.0
C TEXT$22_0/m2_13680_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$1_0/m1_4800_0# TEXT$23_0/m1_7200_0# 0.0
C TEXT$4_0/m3_12000_0# TEXT$22_0/m2_15120_0# 0.0
C TEXT$22_0/m2_5760_0# TEXT$23_0/m1_5760_0# 0.4
C TEXT$23_0/m1_17280_0# TEXT$20_0/m3_17280_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$21_0/m4_7920_720# 0.0
C TEXT$8_0/m4_0_0# TEXT$8_0/m4_960_0# 0.2
C TEXT$23_0/m1_14400_0# TEXT$22_0/m2_14400_0# 0.4
C TEXT$4_0/m3_0_0# TEXT$22_0/m2_2160_0# 0.0
C TEXT$24_0/m3_9600_0# TEXT$7_0/m2_10560_0# 0.0
C TEXT$24_0/m3_10560_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$8_0/m4_6720_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$6_0/m4_3600_0# 0.0
C TEXT$24_0/m3_5760_0# TEXT$23_0/m1_9360_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$6_0/m4_3600_0# 0.0
C TEXT$20_0/m3_8640_0# TEXT$7_0/m2_3840_0# 0.0
C TEXT$23_0/m1_15120_0# TEXT$24_0/m3_10560_0# 0.0
C TEXT$1_0/m1_7200_0# TEXT$21_0/m4_10080_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$4_0/m3_6000_0# 0.3
C TEXT$22_0/m2_10080_0# TEXT$20_0/m3_10080_0# 0.4
C TEXT$22_0/m2_14400_0# TEXT$21_0/m4_15120_0# 0.0
C TEXT$4_0/m3_10800_0# TEXT$6_0/m4_10800_0# 1.2
C TEXT$20_0/m3_3780_0# TEXT$20_0/m3_4320_0# 0.1
C TEXT$23_0/m1_12960_0# TEXT$6_0/m4_10800_0# 0.0
C TEXT$22_0/m2_3780_0# TEXT$21_0/m4_2880_720# 0.0
C TEXT$22_0/m2_2880_720# TEXT$21_0/m4_3780_0# 0.0
C TEXT$6_0/m4_0_0# TEXT$3_0/m2_0_0# 0.0
C TEXT$23_0/m1_17280_0# TEXT$22_0/m2_16560_0# 0.0
C TEXT$20_0/m3_9360_0# TEXT$23_0/m1_9360_0# 0.0
C TEXT$21_0/m4_2880_720# TEXT$23_0/m1_2160_0# 0.0
C VDD TEXT$8_0/m4_960_0# 0.0
C TEXT$24_0/m3_3840_0# TEXT$7_0/m2_3840_0# 0.7
C TEXT$8_0/m4_960_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$21_0/m4_10080_0# TEXT$9_0/m1_5760_0# 0.0
C TEXT$20_0/m3_6480_0# TEXT$21_0/m4_6480_0# 0.4
C TEXT$1_0/m1_9600_0# TEXT$3_0/m2_9600_0# 1.0
C TEXT$1_0/m1_8400_0# TEXT$1_0/m1_9600_0# 0.3
C TEXT$3_0/m2_9600_0# TEXT$3_0/m2_10800_0# 0.1
C TEXT$22_0/m2_10800_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$4_0/m3_12000_0# TEXT$21_0/m4_14400_0# 0.0
C TEXT$8_0/m4_5760_0# TEXT$24_0/m3_6720_0# 0.0
C TEXT$22_0/m2_9360_0# TEXT$21_0/m4_9360_0# 0.0
C TEXT$20_0/m3_10800_0# TEXT$20_0/m3_11700_0# 0.1
C TEXT$21_0/m4_5760_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$23_0/m1_13680_0# TEXT$21_0/m4_14400_0# 0.0
C TEXT$24_0/m3_4800_960# TEXT$23_0/m1_9360_0# 0.0
C TEXT$24_0/m3_5760_0# TEXT$23_0/m1_10080_0# 0.0
C sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# 0.0
C TEXT$4_0/m3_2400_0# TEXT$3_0/m2_2400_0# 1.0
C TEXT$22_0/m2_4320_0# TEXT$3_0/m2_2400_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$23_0/m1_7200_0# 0.0
C TEXT$20_0/m3_10080_0# TEXT$8_0/m4_5760_0# 0.0
C TEXT$20_0/m3_16560_0# TEXT$22_0/m2_15840_0# 0.0
C TEXT$4_0/m3_0_0# TEXT$21_0/m4_2160_0# 0.0
C TEXT$22_0/m2_2880_720# TEXT$21_0/m4_2880_720# 0.0
C TEXT$21_0/m4_10800_0# TEXT$24_0/m3_6720_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$23_0/m1_7200_0# 0.0
C TEXT$20_0/m3_9360_0# TEXT$23_0/m1_10080_0# 0.0
C TEXT$1_0/m1_6000_0# TEXT$6_0/m4_4800_0# 0.0
C TEXT$8_0/m4_2160_0# TEXT$24_0/m3_960_0# 0.0
C TEXT$8_0/m4_4800_960# TEXT$9_0/m1_4800_960# 0.0
C VDD TEXT$9_0/m1_3840_0# 0.0
C TEXT$4_0/m3_7200_0# TEXT$3_0/m2_7200_0# 0.7
C TEXT$1_0/m1_6000_0# TEXT$4_0/m3_7200_0# 0.0
C TEXT$22_0/m2_7200_0# TEXT$8_0/m4_2880_0# 0.0
C TEXT$20_0/m3_10800_0# TEXT$21_0/m4_10080_0# 0.0
C TEXT$20_0/m3_10080_0# TEXT$21_0/m4_10800_0# 0.0
C TEXT$21_0/m4_7200_0# TEXT$7_0/m2_2880_0# 0.0
C TEXT$24_0/m3_0_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$21_0/m4_2880_720# TEXT$21_0/m4_3780_0# 0.1
C TEXT$20_0/m3_720_0# TEXT$20_0/m3_1440_0# 0.3
C TEXT$1_0/m1_7200_0# TEXT$23_0/m1_9360_0# 0.0
C TEXT$9_0/m1_9600_0# TEXT$7_0/m2_10560_0# 0.0
C TEXT$9_0/m1_10560_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$8_0/m4_2160_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$22_0/m2_11700_0# TEXT$24_0/m3_6720_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$22_0/m2_3780_0# 0.0
C VDD TEXT$8_0/m4_3840_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$20_0/m3_8640_0# 0.1
C VDD TEXT$8_0/m4_7680_0# 0.0
C TEXT$4_0/m3_4800_0# TEXT$20_0/m3_7200_0# 0.0
C TEXT$8_0/m4_2160_0# TEXT$9_0/m1_960_0# 0.0
C TEXT$23_0/m1_15120_0# TEXT$9_0/m1_10560_0# 0.0
C TEXT$3_0/m2_6000_0# TEXT$23_0/m1_7920_720# 0.0
C TEXT$1_0/m1_0_0# TEXT$20_0/m3_2880_720# 0.0
C TEXT$22_0/m2_6480_0# TEXT$20_0/m3_7200_0# 0.0
C TEXT$6_0/m4_3600_0# TEXT$6_0/m4_2400_0# 0.2
C TEXT$4_0/m3_6000_0# TEXT$22_0/m2_8640_0# 0.0
C TEXT$7_0/m2_960_0# TEXT$7_0/m2_2160_0# 0.1
C VDD TEXT$7_0/m2_9600_0# 0.0
C TEXT$24_0/m3_7680_0# TEXT$24_0/m3_6720_0# 0.3
C TEXT$20_0/m3_10800_0# TEXT$22_0/m2_10800_0# 0.4
C TEXT$7_0/m2_5760_0# TEXT$9_0/m1_4800_960# 0.0
C TEXT$20_0/m3_15840_0# TEXT$21_0/m4_15840_0# 0.4
C TEXT$22_0/m2_9360_0# TEXT$22_0/m2_10080_0# 0.1
C TEXT$1_0/m1_3600_0# TEXT$3_0/m2_3600_0# 1.1
C TEXT$21_0/m4_9360_0# TEXT$21_0/m4_10080_0# 0.1
C TEXT$24_0/m3_2880_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$22_0/m2_14400_0# TEXT$7_0/m2_10560_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$24_0/m3_3840_0# 0.0
C VDD TEXT$24_0/m3_2160_0# 0.0
C TEXT$24_0/m3_2160_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$22_0/m2_8640_0# TEXT$23_0/m1_9360_0# 0.0
C TEXT$23_0/m1_18000_0# TEXT$20_0/m3_18000_0# 0.0
C TEXT$24_0/m3_5760_0# TEXT$7_0/m2_4800_960# 0.0
C TEXT$8_0/m4_6720_0# TEXT$8_0/m4_7680_0# 0.3
C TEXT$1_0/m1_7200_0# TEXT$23_0/m1_10080_0# 0.0
C TEXT$23_0/m1_15120_0# TEXT$22_0/m2_15120_0# 0.4
C TEXT$21_0/m4_7200_0# TEXT$23_0/m1_7200_0# 0.0
C TEXT$8_0/m4_7680_0# TEXT$7_0/m2_6720_0# 0.0
C TEXT$4_0/m3_7200_0# TEXT$20_0/m3_10080_0# 0.0
C TEXT$20_0/m3_9360_0# TEXT$7_0/m2_4800_960# 0.0
C TEXT$20_0/m3_2160_0# TEXT$3_0/m2_0_0# 0.0
C TEXT$22_0/m2_7200_0# TEXT$6_0/m4_4800_0# 0.0
C TEXT$1_0/m1_8400_0# TEXT$21_0/m4_10800_0# 0.0
C TEXT$21_0/m4_5760_0# TEXT$24_0/m3_960_0# 0.0
C TEXT$22_0/m2_15120_0# TEXT$21_0/m4_15840_0# 0.0
C TEXT$4_0/m3_6000_0# TEXT$22_0/m2_7920_720# 0.0
C TEXT$20_0/m3_4320_0# TEXT$20_0/m3_5760_0# 0.0
C TEXT$23_0/m1_7920_720# TEXT$9_0/m1_3840_0# 0.0
C TEXT$6_0/m4_1200_0# TEXT$3_0/m2_1200_0# 0.0
C TEXT$4_0/m3_1200_0# TEXT$21_0/m4_3780_0# 0.0
C TEXT$23_0/m1_10080_0# TEXT$9_0/m1_5760_0# 0.0
C TEXT$23_0/m1_13680_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$4_0/m3_12000_0# TEXT$23_0/m1_15120_0# 0.0
C TEXT$1_0/m1_6000_0# TEXT$20_0/m3_7920_720# 0.0
C TEXT$24_0/m3_4800_960# TEXT$7_0/m2_4800_960# 0.4
C TEXT$20_0/m3_15120_0# TEXT$8_0/m4_10560_0# 0.0
C TEXT$20_0/m3_7200_0# TEXT$21_0/m4_7200_0# 0.4
C TEXT$1_0/m1_9600_0# TEXT$1_0/m1_10800_0# 0.1
C TEXT$21_0/m4_14400_0# TEXT$7_0/m2_9600_0# 0.0
C TEXT$1_0/m1_8400_0# TEXT$22_0/m2_11700_0# 0.0
C TEXT$1_0/m1_10800_0# TEXT$3_0/m2_10800_0# 1.2
C TEXT$3_0/m2_10800_0# TEXT$3_0/m2_12000_0# 0.1
C TEXT$9_0/m1_5760_0# TEXT$9_0/m1_6720_0# 0.2
C TEXT$22_0/m2_11700_0# TEXT$3_0/m2_9600_0# 0.0
C TEXT$21_0/m4_5760_0# TEXT$9_0/m1_960_0# 0.0
C TEXT$21_0/m4_8640_0# TEXT$7_0/m2_3840_0# 0.0
C TEXT$23_0/m1_8640_0# TEXT$7_0/m2_3840_0# 0.0
C TEXT$22_0/m2_10080_0# TEXT$21_0/m4_10080_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$20_0/m3_12960_0# 0.0
C TEXT$23_0/m1_14400_0# TEXT$21_0/m4_15120_0# 0.0
C TEXT$4_0/m3_3600_0# TEXT$3_0/m2_3600_0# 1.1
C TEXT$22_0/m2_5760_0# TEXT$3_0/m2_3600_0# 0.0
C TEXT$20_0/m3_17280_0# TEXT$22_0/m2_16560_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$23_0/m1_7200_0# 0.0
C TEXT$1_0/m1_1200_0# TEXT$20_0/m3_4320_0# 0.0
C TEXT$22_0/m2_4320_0# TEXT$24_0/m3_0_0# 0.0
C TEXT$1_0/m1_7200_0# TEXT$6_0/m4_6000_0# 0.0
C TEXT$6_0/m4_7200_0# TEXT$3_0/m2_7200_0# 0.0
C TEXT$7_0/m2_0_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$22_0/m2_17280_0# TEXT$23_0/m1_17280_0# 0.4
C TEXT$1_0/m1_7200_0# TEXT$4_0/m3_8400_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$3_0/m2_8400_0# 1.1
C TEXT$6_0/m4_4800_0# TEXT$21_0/m4_7920_720# 0.0
C TEXT$22_0/m2_10080_0# TEXT$22_0/m2_10800_0# 0.2
C TEXT$20_0/m3_11700_0# TEXT$21_0/m4_10800_0# 0.0
C TEXT$8_0/m4_4800_960# TEXT$24_0/m3_5760_0# 0.0
C TEXT$20_0/m3_10800_0# TEXT$9_0/m1_6720_0# 0.0
C TEXT$7_0/m2_960_0# TEXT$23_0/m1_5760_0# 0.0
C TEXT$20_0/m3_720_0# TEXT$22_0/m2_0_0# 0.0
C TEXT$1_0/m1_2400_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$24_0/m3_2160_0# TEXT$8_0/m4_960_0# 0.0
C TEXT$1_0/m1_0_0# TEXT$23_0/m1_2880_720# 0.0
C VDD PD 0.2
C TEXT$21_0/m4_11700_0# TEXT$3_0/m2_8400_0# 0.0
C TEXT$21_0/m4_10080_0# TEXT$8_0/m4_5760_0# 0.0
C TEXT$20_0/m3_9360_0# TEXT$8_0/m4_4800_960# 0.0
C TEXT$7_0/m2_4800_960# TEXT$9_0/m1_5760_0# 0.0
C TEXT$8_0/m4_3840_0# TEXT$9_0/m1_3840_0# 0.0
C TEXT$22_0/m2_6480_0# TEXT$23_0/m1_6480_0# 0.4
C TEXT$8_0/m4_2160_0# TEXT$9_0/m1_2880_0# 0.0
C TEXT$6_0/m4_0_0# TEXT$22_0/m2_2160_0# 0.0
C TEXT$22_0/m2_8640_0# TEXT$6_0/m4_6000_0# 0.0
C TEXT$8_0/m4_9600_0# TEXT$8_0/m4_10560_0# 0.2
C TEXT$22_0/m2_7920_720# TEXT$20_0/m3_7200_0# 0.0
C TEXT$22_0/m2_7200_0# TEXT$20_0/m3_7920_720# 0.0
C TEXT$20_0/m3_3780_0# TEXT$3_0/m2_1200_0# 0.0
C TEXT$4_0/m3_7200_0# TEXT$22_0/m2_9360_0# 0.0
C TEXT$7_0/m2_2160_0# TEXT$7_0/m2_2880_0# 0.1
C TEXT$22_0/m2_8640_0# TEXT$7_0/m2_4800_960# 0.0
C TEXT$1_0/m1_10800_0# TEXT$20_0/m3_12960_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$22_0/m2_11700_0# 0.2
C TEXT$1_0/m1_0_0# TEXT$1_0/m1_1200_0# 0.2
C TEXT$20_0/m3_16560_0# TEXT$21_0/m4_16560_0# 0.4
C TEXT$1_0/m1_4800_0# TEXT$3_0/m2_4800_0# 1.1
C TEXT$21_0/m4_10080_0# TEXT$21_0/m4_10800_0# 0.2
C TEXT$3_0/m2_8400_0# TEXT$23_0/m1_10800_0# 0.0
C TEXT$8_0/m4_4800_960# TEXT$24_0/m3_4800_960# 0.4
C VDD TEXT$24_0/m3_3840_0# 0.0
C TEXT$24_0/m3_5760_0# TEXT$7_0/m2_5760_0# 0.7
C TEXT$24_0/m3_2880_0# TEXT$9_0/m1_2880_0# 0.0
C TEXT$22_0/m2_10080_0# TEXT$23_0/m1_9360_0# 0.0
C TEXT$20_0/m3_11700_0# TEXT$24_0/m3_7680_0# 0.0
C TEXT$21_0/m4_6480_0# TEXT$3_0/m2_3600_0# 0.0
C TEXT$3_0/m2_10800_0# TEXT$6_0/m4_12000_0# 0.0
C TEXT$23_0/m1_11700_0# TEXT$24_0/m3_6720_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$21_0/m4_8640_0# 0.0
C TEXT$20_0/m3_10080_0# TEXT$6_0/m4_7200_0# 0.0
C TEXT$4_0/m3_8400_0# TEXT$20_0/m3_10800_0# 0.0
C TEXT$22_0/m2_7920_720# TEXT$6_0/m4_6000_0# 0.0
C TEXT$22_0/m2_10800_0# TEXT$21_0/m4_10800_0# 0.0
C TEXT$20_0/m3_0_0# TEXT$21_0/m4_720_0# 0.0
C TEXT$22_0/m2_15840_0# TEXT$21_0/m4_16560_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$20_0/m3_6480_0# 0.2
C TEXT$1_0/m1_0_0# TEXT$3_0/m2_0_0# 1.1
C TEXT$4_0/m3_2400_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$6_0/m4_2400_0# TEXT$3_0/m2_2400_0# 0.0
C M_0/a_404041_244568# VDD 1.7
C TEXT$23_0/m1_14400_0# TEXT$7_0/m2_10560_0# 0.0
C TEXT$20_0/m3_4320_0# TEXT$23_0/m1_4320_0# 0.0
C TEXT$22_0/m2_4320_0# TEXT$21_0/m4_4320_0# 0.0
C TEXT$20_0/m3_10800_0# TEXT$21_0/m4_11700_0# 0.0
C TEXT$24_0/m3_9600_0# TEXT$8_0/m4_10560_0# 0.0
C TEXT$6_0/m4_0_0# TEXT$21_0/m4_2160_0# 0.0
C TEXT$22_0/m2_10080_0# TEXT$23_0/m1_10080_0# 0.4
C TEXT$24_0/m3_960_0# TEXT$7_0/m2_0_0# 0.0
C TEXT$8_0/m4_2880_0# TEXT$7_0/m2_2880_0# 0.0
C TEXT$21_0/m4_7200_0# TEXT$23_0/m1_6480_0# 0.0
C TEXT$20_0/m3_5760_0# TEXT$23_0/m1_5760_0# 0.0
C TEXT$20_0/m3_7920_720# TEXT$21_0/m4_7920_720# 0.2
C TEXT$1_0/m1_10800_0# TEXT$1_0/m1_12000_0# 0.1
C TEXT$21_0/m4_15120_0# TEXT$7_0/m2_10560_0# 0.0
C TEXT$1_0/m1_12000_0# TEXT$3_0/m2_12000_0# 1.1
C TEXT$4_0/m3_7200_0# TEXT$21_0/m4_10080_0# 0.0
C TEXT$22_0/m2_12960_0# TEXT$3_0/m2_10800_0# 0.0
C TEXT$22_0/m2_10800_0# TEXT$22_0/m2_11700_0# 0.1
C TEXT$21_0/m4_6480_0# TEXT$9_0/m1_2160_0# 0.0
C TEXT$21_0/m4_9360_0# TEXT$7_0/m2_4800_960# 0.0
C TEXT$20_0/m3_12960_0# TEXT$20_0/m3_13680_0# 0.2
C PD0 2.4
R PD 22
= PD via_dev_0/m1_0_0#
= PD sc_tieh_tiel$1_0/tieH
= PD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/Z
= PD via_dev$42_0/m2_0_0#
= PD m2_516942_218066#
C VBIAS0 21.4
R VBIAS 578
C VIN0 21.6
R VIN 578
C VCM_OUT0 90.4
R VCM_OUT 135
= VCM_OUT via_dev$35_2/m2_0_0#
= VCM_OUT m4_420113_244057#
= VCM_OUT via_dev$34_0/m2_0_0#
= VCM_OUT M_0/a_411044_242557#
C BCM_OUT0 83.5
R BCM_OUT 135
= BCM_OUT via_dev$35_3/m2_0_0#
= BCM_OUT m4_420120_253237#
= BCM_OUT via_dev$34_1/m2_0_0#
= BCM_OUT M_0/a_411044_251737#
C CCM_OUT0 77.4
R CCM_OUT 192
= CCM_OUT via_dev$35_5/m2_0_0#
= CCM_OUT m4_420104_257713#
= CCM_OUT via_dev$34_2/m2_0_0#
= CCM_OUT M_0/a_409818_256643#
C VIN_OUT0 75.9
R VIN_OUT 223
= VIN_OUT via_dev$35_4/m2_0_0#
= VIN_OUT m4_420119_263354#
= VIN_OUT via_dev$34_3/m2_0_0#
= VIN_OUT M_0/a_404831_244568#
R a_510132_239389# 1400
R a_510063_259404# 1400
C TEXT$1_0/m1_12000_0#0 1.7
C TEXT$1_0/m1_10800_0#0 1.6
C TEXT$1_0/m1_9600_0#0 1.5
C TEXT$1_0/m1_8400_0#0 1.6
C TEXT$1_0/m1_7200_0#0 1.0
C TEXT$1_0/m1_6000_0#0 1.5
C TEXT$1_0/m1_4800_0#0 1.4
C TEXT$1_0/m1_3600_0#0 1.5
C TEXT$1_0/m1_2400_0#0 1.4
C TEXT$1_0/m1_1200_0#0 1.5
C TEXT$1_0/m1_0_0#0 1.6
C M_0/a_410724_251737#0 2.9
R M_0/a_410724_251737# 107
C M_0/a_410134_251737#0 6.4
R M_0/a_410134_251737# 219
C M_0/a_409498_256643#0 8.5
R M_0/a_409498_256643# 340
C M_0/a_409618_260539#0 8.4
R M_0/a_409618_260539# 335
C M_0/a_404041_244568#0 14.1
R M_0/a_404041_244568# 489
C M_0/a_403251_244568#0 5.1
R M_0/a_403251_244568# 293
C M_0/a_402461_244568#0 8.1
R M_0/a_402461_244568# 292
C a_498947_268180#0 209.0
R a_498947_268180# 881
= a_498947_268180# via_dev$35_6/m2_0_0#
= a_498947_268180# m4_399395_244477#
= a_498947_268180# via_dev$35_7/m2_0_0#
= a_498947_268180# m2_399395_243478#
= a_498947_268180# M_0/a_401271_243528#
C M_0/a_404311_244568#0 0.2
R M_0/a_404311_244568# 272
C M_0/a_403521_244568#0 0.0
R M_0/a_403521_244568# 272
C M_0/a_402731_244568#0 0.0
R M_0/a_402731_244568# 272
C M_0/a_401941_244568#0 0.0
R M_0/a_401941_244568# 272
C M_0/a_401151_244568#0 2.6
R M_0/a_401151_244568# 1220
C m4_400150_261569#0 16.5
R m4_400150_261569# 601
= m4_400150_261569# via_dev$35_1/m2_0_0#
= m4_400150_261569# M_0/a_409618_256263#
= m4_400150_261569# via_dev$35_0/m2_0_0#
= m4_400150_261569# m2_397020_261569#
= m4_400150_261569# M_0/a_395682_259299#
C M_0/a_395162_259299#0 0.3
R M_0/a_395162_259299# 260
C M_0/a_383940_262205#0 4.9
R M_0/a_383940_262205# 2090
C M_0/a_383620_262205#0 2.8
R M_0/a_383620_262205# 191
C M_0/a_377450_262205#0 40.1
R M_0/a_377450_262205# 2962
C M_0/a_374398_259299#0 12.9
R M_0/a_374398_259299# 2054
C a_499016_248165#0 232.3
R a_499016_248165# 2377
= a_499016_248165# via_dev$32_1/m2_0_0#
= a_499016_248165# m3_420393_272672#
= a_499016_248165# M_0/a_365828_259091#
C M_0/a_373878_259299#0 0.2
R M_0/a_373878_259299# 260
C M_0/a_386992_259299#0 3.2
R M_0/a_386992_259299# 3505
C M_0/a_365708_259299#0 3.2
R M_0/a_365708_259299# 3505
C TEXT$3_0/m2_12000_0#0 1.1
C TEXT$3_0/m2_10800_0#0 1.0
C TEXT$3_0/m2_9600_0#0 0.9
C TEXT$3_0/m2_8400_0#0 1.0
C TEXT$3_0/m2_7200_0#0 0.7
C TEXT$3_0/m2_6000_0#0 0.9
C TEXT$3_0/m2_4800_0#0 0.8
C TEXT$3_0/m2_3600_0#0 0.9
C TEXT$3_0/m2_2400_0#0 0.9
C TEXT$3_0/m2_1200_0#0 0.9
C TEXT$3_0/m2_0_0#0 1.0
C TEXT$21_0/m4_18000_0#0 0.4
C TEXT$21_0/m4_17280_0#0 0.3
C TEXT$21_0/m4_16560_0#0 0.3
C TEXT$21_0/m4_15840_0#0 0.3
C TEXT$21_0/m4_15120_0#0 0.3
C TEXT$21_0/m4_14400_0#0 0.3
C TEXT$21_0/m4_13680_0#0 0.3
C TEXT$21_0/m4_12960_0#0 0.3
C TEXT$21_0/m4_11700_0#0 0.2
C TEXT$21_0/m4_10800_0#0 0.3
C TEXT$21_0/m4_10080_0#0 0.3
C TEXT$21_0/m4_9360_0#0 0.3
C TEXT$21_0/m4_8640_0#0 0.3
C TEXT$21_0/m4_7920_720#0 0.2
C TEXT$21_0/m4_7200_0#0 0.3
C TEXT$21_0/m4_6480_0#0 0.3
C TEXT$21_0/m4_5760_0#0 0.3
C TEXT$21_0/m4_4320_0#0 0.3
C TEXT$21_0/m4_3780_0#0 0.2
C TEXT$21_0/m4_2880_720#0 0.2
C TEXT$21_0/m4_2160_0#0 0.3
C TEXT$21_0/m4_1440_0#0 0.3
C TEXT$21_0/m4_720_0#0 0.3
C TEXT$21_0/m4_0_0#0 0.4
C TEXT$23_0/m1_18000_0#0 0.7
C TEXT$23_0/m1_17280_0#0 0.7
C TEXT$23_0/m1_16560_0#0 0.6
C TEXT$23_0/m1_15840_0#0 0.7
C TEXT$23_0/m1_15120_0#0 0.6
C TEXT$23_0/m1_14400_0#0 0.7
C TEXT$23_0/m1_13680_0#0 0.6
C TEXT$23_0/m1_12960_0#0 0.7
C TEXT$23_0/m1_11700_0#0 0.4
C TEXT$23_0/m1_10800_0#0 0.7
C TEXT$23_0/m1_10080_0#0 0.7
C TEXT$23_0/m1_9360_0#0 0.7
C TEXT$23_0/m1_8640_0#0 0.7
C TEXT$23_0/m1_7920_720#0 0.5
C TEXT$23_0/m1_7200_0#0 0.6
C TEXT$23_0/m1_6480_0#0 0.7
C TEXT$23_0/m1_5760_0#0 0.7
C TEXT$23_0/m1_4320_0#0 0.7
C TEXT$23_0/m1_3780_0#0 0.4
C TEXT$23_0/m1_2880_720#0 0.5
C TEXT$23_0/m1_2160_0#0 0.7
C TEXT$23_0/m1_1440_0#0 0.7
C TEXT$23_0/m1_720_0#0 0.6
C TEXT$23_0/m1_0_0#0 0.8
C m3_419992_265695#0 234.5
R m3_419992_265695# 783
= m3_419992_265695# via_dev$32_0/m2_0_0#
= m3_419992_265695# m2_477527_223220#
= m3_419992_265695# via_dev$33_0/m2_0_0#
= m3_419992_265695# M_0/a_365828_265695#
= m3_419992_265695# io_secondary_5p0$1_0/m1_499212_228525#
= m3_419992_265695# io_secondary_5p0$1_0/diode_pd2nw_06v0_5DG9HC_0/a_507479_219793#
= m3_419992_265695# io_secondary_5p0$1_0/diode_pd2nw_06v0_5DG9HC_0/a_505263_219793#
= m3_419992_265695# io_secondary_5p0$1_0/diode_pd2nw_06v0_5DG9HC_0/a_503047_219793#
= m3_419992_265695# io_secondary_5p0$1_0/diode_pd2nw_06v0_5DG9HC_0/a_500831_219793#
= m3_419992_265695# io_secondary_5p0$1_0/ppolyf_u_9H3LNU_0/a_n224793_504053#
= m3_419992_265695# io_secondary_5p0$1_0/diode_nd2ps_06v0_MV3SZ3_0/a_507503_219793#
= m3_419992_265695# io_secondary_5p0$1_0/diode_nd2ps_06v0_MV3SZ3_0/a_505271_219793#
= m3_419992_265695# io_secondary_5p0$1_0/diode_nd2ps_06v0_MV3SZ3_0/a_503039_219793#
= m3_419992_265695# io_secondary_5p0$1_0/diode_nd2ps_06v0_MV3SZ3_0/a_500807_219793#
R io_secondary_5p0$1_0/ppolyf_u_9H3LNU_0/a_n224793_504155# 1400
C EN0 6.2
R EN 584
= EN io_secondary_5p0$1_0/m1_512035_219553#
= EN io_secondary_5p0$1_0/ppolyf_u_9H3LNU_0/a_n224793_506155#
C TEXT$7_0/m2_10560_0#0 0.8
C TEXT$7_0/m2_9600_0#0 0.7
C TEXT$7_0/m2_7680_0#0 0.7
C TEXT$7_0/m2_6720_0#0 0.7
C TEXT$7_0/m2_5760_0#0 0.7
C TEXT$7_0/m2_4800_960#0 0.5
C TEXT$7_0/m2_3840_0#0 0.7
C TEXT$7_0/m2_2880_0#0 0.6
C TEXT$7_0/m2_2160_0#0 0.4
C TEXT$7_0/m2_960_0#0 0.7
C TEXT$7_0/m2_0_0#0 0.7
C TEXT$9_0/m1_10560_0#0 1.2
C TEXT$9_0/m1_9600_0#0 1.1
C TEXT$9_0/m1_7680_0#0 1.1
C TEXT$9_0/m1_6720_0#0 1.1
C TEXT$9_0/m1_5760_0#0 1.0
C TEXT$9_0/m1_4800_960#0 0.8
C TEXT$9_0/m1_3840_0#0 1.1
C TEXT$9_0/m1_2880_0#0 1.0
C TEXT$9_0/m1_2160_0#0 0.6
C TEXT$9_0/m1_960_0#0 1.1
C TEXT$9_0/m1_0_0#0 1.1
R TEXT$9_0/VSUBS 72427
= TEXT$9_0/VSUBS DNWell_Rect_0/w_407433_240888#
= TEXT$9_0/VSUBS w_407433_240888#
= TEXT$9_0/VSUBS via_dev$35_4/VSUBS
= TEXT$9_0/VSUBS via_dev$34_3/VSUBS
= TEXT$9_0/VSUBS via_dev$35_1/VSUBS
= TEXT$9_0/VSUBS via_dev$35_0/VSUBS
= TEXT$9_0/VSUBS via_dev$35_5/VSUBS
= TEXT$9_0/VSUBS via_dev$34_2/VSUBS
= TEXT$9_0/VSUBS via_dev$37_2/VSUBS
= TEXT$9_0/VSUBS via_dev$37_2/m1_0_0#
= TEXT$9_0/VSUBS via_dev$35_3/VSUBS
= TEXT$9_0/VSUBS via_dev$34_1/VSUBS
= TEXT$9_0/VSUBS via_dev$41_1/VSUBS
= TEXT$9_0/VSUBS via_dev$35_7/VSUBS
= TEXT$9_0/VSUBS via_dev$35_2/VSUBS
= TEXT$9_0/VSUBS via_dev$34_0/VSUBS
= TEXT$9_0/VSUBS M_0/a_376520_259212#
= TEXT$9_0/VSUBS DNWell_Rect_0/a_406361_239816#
= TEXT$9_0/VSUBS via_dev$37_1/VSUBS
= TEXT$9_0/VSUBS via_dev$37_1/m1_0_0#
= TEXT$9_0/VSUBS via_dev$45_0/m1_0_0#
= TEXT$9_0/VSUBS m2_514376_217140#
= TEXT$9_0/VSUBS via_dev$37_0/m1_0_0#
= TEXT$9_0/VSUBS m1_507881_217140#
= TEXT$9_0/VSUBS m3_410146_285414#
= TEXT$9_0/VSUBS via_dev$41_0/VSUBS
= TEXT$9_0/VSUBS via_dev_0/VSUBS
= TEXT$9_0/VSUBS via_dev$44_0/VSUBS
= TEXT$9_0/VSUBS sc_tieh_tiel_0/VSUBS
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/VSS
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/VPW
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/VSS
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/VPW
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/VSS
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__filltie$1_1/VSS
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__filltie$1_0/VSS
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/via_dev$43_1/VSUBS
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/via_dev$43_0/VSUBS
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/VSUBS
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/via_dev$43_1/m1_0_0#
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/m1_396908_517398#
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/via_dev$43_0/m1_0_0#
= TEXT$9_0/VSUBS sc_tieh_tiel$1_0/m2_396908_515382#
= TEXT$9_0/VSUBS via_dev$42_0/VSUBS
= TEXT$9_0/VSUBS via_dev$45_0/VSUBS
= TEXT$9_0/VSUBS TEXT$6_0/VSUBS
= TEXT$9_0/VSUBS TEXT$4_0/VSUBS
= TEXT$9_0/VSUBS TEXT$3_0/VSUBS
= TEXT$9_0/VSUBS TEXT$1_0/VSUBS
= TEXT$9_0/VSUBS via_dev$37_0/VSUBS
= TEXT$9_0/VSUBS io_secondary_5p0$1_0/VSUBS
= TEXT$9_0/VSUBS io_secondary_5p0$1_0/diode_pd2nw_06v0_5DG9HC_0/a_500511_219473#
= TEXT$9_0/VSUBS io_secondary_5p0$1_0/ppolyf_u_9H3LNU_0/VSUBS
= TEXT$9_0/VSUBS io_secondary_5p0$1_0/diode_nd2ps_06v0_MV3SZ3_0/a_500655_219641#
= TEXT$9_0/VSUBS io_secondary_5p0$1_0/m1_497955_215963#
= TEXT$9_0/VSUBS TEXT$21_0/VSUBS
= TEXT$9_0/VSUBS TEXT$20_0/VSUBS
= TEXT$9_0/VSUBS TEXT$22_0/VSUBS
= TEXT$9_0/VSUBS TEXT$23_0/VSUBS
= TEXT$9_0/VSUBS TEXT$8_0/VSUBS
= TEXT$9_0/VSUBS TEXT$24_0/VSUBS
= TEXT$9_0/VSUBS TEXT$7_0/VSUBS
= TEXT$9_0/VSUBS a_344599_211617#
C TEXT$20_0/m3_18000_0#0 0.4
C TEXT$20_0/m3_17280_0#0 0.3
C TEXT$20_0/m3_16560_0#0 0.3
C TEXT$20_0/m3_15840_0#0 0.3
C TEXT$20_0/m3_15120_0#0 0.3
C TEXT$20_0/m3_14400_0#0 0.3
C TEXT$20_0/m3_13680_0#0 0.3
C TEXT$20_0/m3_12960_0#0 0.4
C TEXT$20_0/m3_11700_0#0 0.2
C TEXT$20_0/m3_10800_0#0 0.3
C TEXT$20_0/m3_10080_0#0 0.3
C TEXT$20_0/m3_9360_0#0 0.3
C TEXT$20_0/m3_8640_0#0 0.3
C TEXT$20_0/m3_7920_720#0 0.3
C TEXT$20_0/m3_7200_0#0 0.3
C TEXT$20_0/m3_6480_0#0 0.3
C TEXT$20_0/m3_5760_0#0 0.4
C TEXT$20_0/m3_4320_0#0 0.4
C TEXT$20_0/m3_3780_0#0 0.2
C TEXT$20_0/m3_2880_720#0 0.3
C TEXT$20_0/m3_2160_0#0 0.3
C TEXT$20_0/m3_1440_0#0 0.3
C TEXT$20_0/m3_720_0#0 0.3
C TEXT$20_0/m3_0_0#0 0.4
C TEXT$4_0/m3_12000_0#0 0.9
C TEXT$4_0/m3_10800_0#0 0.7
C TEXT$4_0/m3_9600_0#0 0.7
C TEXT$4_0/m3_8400_0#0 0.8
C TEXT$4_0/m3_7200_0#0 0.5
C TEXT$4_0/m3_6000_0#0 0.7
C TEXT$4_0/m3_4800_0#0 0.6
C TEXT$4_0/m3_3600_0#0 0.7
C TEXT$4_0/m3_2400_0#0 0.7
C TEXT$4_0/m3_1200_0#0 0.7
C TEXT$4_0/m3_0_0#0 0.8
C TEXT$22_0/m2_18000_0#0 0.5
C TEXT$22_0/m2_17280_0#0 0.4
C TEXT$22_0/m2_16560_0#0 0.4
C TEXT$22_0/m2_15840_0#0 0.4
C TEXT$22_0/m2_15120_0#0 0.4
C TEXT$22_0/m2_14400_0#0 0.4
C TEXT$22_0/m2_13680_0#0 0.4
C TEXT$22_0/m2_12960_0#0 0.5
C TEXT$22_0/m2_11700_0#0 0.3
C TEXT$22_0/m2_10800_0#0 0.4
C TEXT$22_0/m2_10080_0#0 0.4
C TEXT$22_0/m2_9360_0#0 0.4
C TEXT$22_0/m2_8640_0#0 0.4
C TEXT$22_0/m2_7920_720#0 0.4
C TEXT$22_0/m2_7200_0#0 0.4
C TEXT$22_0/m2_6480_0#0 0.4
C TEXT$22_0/m2_5760_0#0 0.5
C TEXT$22_0/m2_4320_0#0 0.5
C TEXT$22_0/m2_3780_0#0 0.3
C TEXT$22_0/m2_2880_720#0 0.4
C TEXT$22_0/m2_2160_0#0 0.4
C TEXT$22_0/m2_1440_0#0 0.4
C TEXT$22_0/m2_720_0#0 0.4
C TEXT$22_0/m2_0_0#0 0.5
C TEXT$6_0/m4_12000_0#0 0.8
C TEXT$6_0/m4_10800_0#0 0.6
C TEXT$6_0/m4_9600_0#0 0.6
C TEXT$6_0/m4_8400_0#0 0.7
C TEXT$6_0/m4_7200_0#0 0.5
C TEXT$6_0/m4_6000_0#0 0.6
C TEXT$6_0/m4_4800_0#0 0.5
C TEXT$6_0/m4_3600_0#0 0.6
C TEXT$6_0/m4_2400_0#0 0.5
C TEXT$6_0/m4_1200_0#0 0.6
C TEXT$6_0/m4_0_0#0 0.7
C TEXT$24_0/m3_10560_0#0 0.7
C TEXT$24_0/m3_9600_0#0 0.6
C TEXT$24_0/m3_7680_0#0 0.5
C TEXT$24_0/m3_6720_0#0 0.5
C TEXT$24_0/m3_5760_0#0 0.5
C TEXT$24_0/m3_4800_960#0 0.4
C TEXT$24_0/m3_3840_0#0 0.6
C TEXT$24_0/m3_2880_0#0 0.5
C TEXT$24_0/m3_2160_0#0 0.3
C TEXT$24_0/m3_960_0#0 0.5
C TEXT$24_0/m3_0_0#0 0.6
C TEXT$8_0/m4_10560_0#0 0.6
C TEXT$8_0/m4_9600_0#0 0.5
C TEXT$8_0/m4_7680_0#0 0.5
C TEXT$8_0/m4_6720_0#0 0.5
C TEXT$8_0/m4_5760_0#0 0.4
C TEXT$8_0/m4_4800_960#0 0.4
C TEXT$8_0/m4_3840_0#0 0.5
C TEXT$8_0/m4_2880_0#0 0.4
C TEXT$8_0/m4_2160_0#0 0.2
C TEXT$8_0/m4_960_0#0 0.4
C TEXT$8_0/m4_0_0#0 0.5
C VDD0 2432.8
R VDD 555999
= VDD via_dev$39_0/m2_0_0#
= VDD via_dev$15_0/m2_0_0#
= VDD via_dev$29_0/m1_0_0#
= VDD m4_409998_292651#
= VDD M_0/w_364522_258756#
= VDD w_345212_212189#
= VDD sc_tieh_tiel$1_0/VDD
= VDD via_dev$41_2/m1_0_0#
= VDD w_498771_268004#
= VDD via_dev$41_1/m1_0_0#
= VDD w_498840_247989#
= VDD via_dev$41_0/m1_0_0#
= VDD m3_510297_218284#
= VDD io_secondary_5p0$1_0/m1_497955_232243#
= VDD io_secondary_5p0$1_0/diode_pd2nw_06v0_5DG9HC_0/w_500655_219617#
= VDD io_secondary_5p0$1_0/ppolyf_u_9H3LNU_0/w_n225009_503837#
= VDD m1_512118_230975#
= VDD sc_tieh_tiel_0/m1_514121_226826#
= VDD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/VDD
= VDD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/VNW
= VDD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/VDD
= VDD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/VNW
= VDD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__filltie$1_1/VDD
= VDD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__filltie$1_0/VDD
C PU0 6.0
R PU 28
= PU via_dev$44_0/m1_0_0#
= PU sc_tieh_tiel$1_0/tieL
= PU sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/ZN
C sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157#0 0.4
R sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# 61
C sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157#0 0.5
R sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# 72
= VSS via_dev$39_0/VSUBS
= VSS via_dev$15_0/VSUBS
= VSS via_dev$29_0/VSUBS
= VSS via_dev$14_0/VSUBS
= VSS via_dev$14_0/m2_0_0#
= VSS via_dev$11_0/VSUBS
= VSS via_dev$11_0/m1_0_0#
= VSS via_dev$36_0/VSUBS
= VSS via_dev$36_0/m1_0_0#
= VSS via_dev$38_0/VSUBS
= VSS via_dev$41_2/VSUBS
= VSS via_dev$38_0/m2_0_0#
= VSS via_dev$35_6/VSUBS
= VSS via_dev$32_1/VSUBS
= VSS via_dev$33_0/VSUBS
= VSS via_dev$32_0/VSUBS
