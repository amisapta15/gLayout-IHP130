* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VIN VSS VDD VOUT_RCCM VOUT_SBCM VOUT_VCM VAUX EN
X0 VAUX a_5777_8307# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X1 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X2 VAUX a_5777_8307# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X3 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0.17441n ps=0.65676m w=4u l=1u
X4 VAUX a_5657_4411# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X5 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X6 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X7 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X8 a_n40012_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X9 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X10 VAUX a_5657_4411# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X11 a_n715_n5930# a_n1505_n5930# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X12 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0.1116n ps=0.40232m w=10u l=2u
X13 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X14 a_n30270_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X15 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X16 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X17 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X18 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X19 a_n195_n5930# VIN a_n715_n5930# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X20 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X21 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X22 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X23 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X24 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X25 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X26 a_75_n5930# a_n1505_n5930# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X27 a_595_n5930# a_595_n5930# a_6293_483# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X28 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X29 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X30 a_1385_n5930# VAUX a_5777_8307# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X31 a_1385_n5930# VAUX a_5777_8307# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X32 a_595_n5930# VIN a_75_n5930# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X33 a_n1505_n5930# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X34 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X35 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X36 a_n29950_3049# a_n39492_5979# a_n30270_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X37 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X38 a_6883_483# a_6293_483# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X39 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X40 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0.27118n ps=0.97416m w=10u l=2u
X41 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X42 a_5777_8307# a_1385_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X43 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X44 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X45 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X46 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X47 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.7971p pd=21.15u as=0 ps=0 w=9.995u l=2u
X48 a_5777_8307# a_1385_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X49 a_n18208_5979# a_n29950_3049# a_n18728_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X50 VOUT_VCM a_n195_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X51 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X52 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X53 VOUT_SBCM a_595_n5930# a_6883_483# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X54 VSS VSS VSS VSS nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X55 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X56 a_n26898_5979# a_n48062_12376# a_n26898_12584# w_n49368_5436# pfet_03v3 ad=5.997p pd=21.19u as=5.997p ps=21.19u w=9.995u l=2u
X57 VSS VSS VSS VSS nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X58 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X59 a_n48182_5979# a_n48062_12376# a_n48182_12584# w_n49368_5436# pfet_03v3 ad=5.997p pd=21.19u as=5.997p ps=21.19u w=9.995u l=2u
X60 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X61 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X62 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X63 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X64 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X65 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X66 a_5657_4411# a_1385_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X67 a_5657_4411# a_1385_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X68 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X69 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X70 VSS VSS VSS VSS nfet_03v3 ad=4.6429p pd=17.17u as=0 ps=0 w=8.005u l=1u
X71 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X72 a_n39492_5979# a_n48062_5772# a_n40012_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X73 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X74 a_n1505_n5930# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X75 a_n1505_n5930# a_n1505_n5930# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X76 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X77 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X78 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X79 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X80 a_n39492_5979# a_n31010_3002# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X81 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X82 VIN VIN a_n1505_n5930# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X83 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X84 a_n1505_n5930# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X85 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X86 a_865_n5930# a_n1505_n5930# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X87 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X88 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X89 a_6293_483# a_6293_483# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X90 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X91 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X92 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X93 a_1385_n5930# VIN a_865_n5930# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X94 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X95 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X96 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X97 a_n195_n5930# a_n195_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X98 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X99 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X100 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X101 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X102 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X103 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X104 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X105 a_n18728_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X106 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.7971p pd=21.15u as=0 ps=0 w=9.995u l=2u
X107 VOUT_RCCM VAUX a_5657_4411# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X108 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X109 VSS VSS VSS VSS nfet_03v3 ad=4.6429p pd=17.17u as=0 ps=0 w=8.005u l=1u
X110 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X111 VOUT_RCCM VAUX a_5657_4411# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X112 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X113 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.7971p pd=21.15u as=0 ps=0 w=9.995u l=2u
X114 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X115 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.7971p pd=21.15u as=0 ps=0 w=9.995u l=2u
X116 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X117 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X118 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X119 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X120 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X121 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X122 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X123 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X124 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X125 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X126 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X127 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X128 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X129 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X130 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
C0 a_1385_n5930# VOUT_RCCM 0.00933f
C1 a_n195_n5930# a_865_n5930# 0.10043f
C2 a_595_n5930# a_865_n5930# 2.02912f
C3 a_n31010_3002# a_n30270_3049# 0.00593f
C4 a_n36440_3049# a_n39492_5979# 36.2174f
C5 a_n48182_5979# a_n39492_5979# 0.06695f
C6 a_595_n5930# VOUT_SBCM 0.2042f
C7 a_1385_n5930# a_75_n5930# 0.13665f
C8 a_595_n5930# a_6293_483# 1.85176f
C9 a_n29950_3049# a_n30270_3049# 1.13457f
C10 w_n49368_5436# a_n48062_5772# 15.1108f
C11 VAUX a_5657_4411# 3.29507f
C12 a_n48062_12376# a_n40012_5979# 0
C13 a_595_n5930# VDD 0.97996f
C14 a_n195_n5930# VDD 1.06408f
C15 VOUT_SBCM a_6293_483# 0.0849f
C16 a_n29950_3049# a_n18208_5979# 0.50367f
C17 a_n195_n5930# a_n1505_n5930# 0.13478f
C18 a_595_n5930# a_n1505_n5930# 0.13836f
C19 a_865_n5930# EN 0.21853f
C20 a_n31010_3002# a_n39492_5979# 0.07262f
C21 a_1385_n5930# a_n715_n5930# 0.13688f
C22 VAUX a_5777_8307# 3.58908f
C23 a_n195_n5930# VIN 0.63325f
C24 a_595_n5930# VIN 0.62256f
C25 a_75_n5930# a_n715_n5930# 0.78447f
C26 a_865_n5930# VDD 5.40929f
C27 a_865_n5930# a_n1505_n5930# 2.19448f
C28 a_n29950_3049# a_n39492_5979# 0.28183f
C29 a_n48182_5979# a_n48062_5772# 29.4854f
C30 a_n26898_5979# a_n29950_3049# 29.5536f
C31 a_n48182_12584# w_n49368_5436# 1.36726f
C32 VIN a_865_n5930# 0.62292f
C33 a_n48182_5979# w_n49368_5436# 47.6849f
C34 a_n39492_5979# a_n40012_5979# 0.85651f
C35 VAUX VOUT_RCCM 0.57679f
C36 a_n18728_5979# a_n29950_3049# 0.99953f
C37 VAUX a_1385_n5930# 1.72199f
C38 EN VDD 7.30305f
C39 EN a_n1505_n5930# 1.62501f
C40 a_n39492_5979# a_n30270_3049# 0.85955f
C41 a_595_n5930# a_6883_483# 1.45997f
C42 a_n26898_5979# a_n48062_12376# 0.70477f
C43 VDD a_n1505_n5930# 31.4897f
C44 a_n26898_12584# a_n48062_12376# 0.5732f
C45 VIN VDD 10.2566f
C46 a_n48182_12584# a_n48182_5979# 0.99741f
C47 VIN a_n1505_n5930# 2.98274f
C48 a_n195_n5930# a_1385_n5930# 0.08093f
C49 a_595_n5930# a_1385_n5930# 0.42594f
C50 a_n26898_5979# a_n18208_5979# 0.06695f
C51 a_n195_n5930# a_75_n5930# 2.03168f
C52 a_595_n5930# a_75_n5930# 2.02098f
C53 VOUT_SBCM a_6883_483# 1.15251f
C54 a_n29950_3049# w_n49368_5436# 15.4156f
C55 a_6883_483# a_6293_483# 0.36588f
C56 a_1385_n5930# a_865_n5930# 1.98101f
C57 a_n40012_5979# a_n48062_5772# 0.99953f
C58 a_n18728_5979# a_n18208_5979# 0.85331f
C59 a_865_n5930# a_75_n5930# 0.74423f
C60 w_n49368_5436# a_n40012_5979# 3.05519f
C61 a_n26898_5979# a_n26898_12584# 0.99741f
C62 a_n26898_5979# a_n18728_5979# 0.98687f
C63 a_n31010_3002# a_n36440_3049# 0.35829f
C64 a_5777_8307# a_5657_4411# 0.36393f
C65 a_n195_n5930# a_n715_n5930# 2.02854f
C66 a_595_n5930# a_n715_n5930# 0.17152f
C67 w_n49368_5436# a_n48062_12376# 5.46416f
C68 EN a_75_n5930# 0.00866f
C69 a_n29950_3049# a_n36440_3049# 0
C70 a_1385_n5930# VDD 2.57265f
C71 a_1385_n5930# a_n1505_n5930# 0.82034f
C72 a_865_n5930# a_n715_n5930# 0.30282f
C73 VOUT_RCCM a_5657_4411# 2.17202f
C74 VDD a_75_n5930# 6.35872f
C75 a_75_n5930# a_n1505_n5930# 1.38044f
C76 a_1385_n5930# VIN 0.55089f
C77 w_n49368_5436# a_n18208_5979# 1.49145f
C78 a_n48182_5979# a_n40012_5979# 0.98687f
C79 a_1385_n5930# a_5657_4411# 0.85546f
C80 VIN a_75_n5930# 0.6318f
C81 a_n39492_5979# a_n48062_5772# 0.50698f
C82 a_n195_n5930# VOUT_VCM 0.20751f
C83 a_n36440_3049# a_n30270_3049# 0.52271f
C84 w_n49368_5436# a_n39492_5979# 1.79624f
C85 a_n26898_5979# w_n49368_5436# 47.7034f
C86 a_n48182_12584# a_n48062_12376# 0.5732f
C87 EN a_n715_n5930# 0.00664f
C88 VOUT_RCCM a_5777_8307# 0.0136f
C89 a_n48182_5979# a_n48062_12376# 0.75535f
C90 w_n49368_5436# a_n26898_12584# 1.375f
C91 a_n31010_3002# a_n29950_3049# 0
C92 a_1385_n5930# a_5777_8307# 3.00275f
C93 a_n18728_5979# w_n49368_5436# 3.05519f
C94 VDD a_n715_n5930# 6.34675f
C95 a_n715_n5930# a_n1505_n5930# 1.68766f
C96 a_595_n5930# a_n195_n5930# 0.53741f
C97 VIN a_n715_n5930# 2.59448f
C98 VOUT_VCM VSS 3.01288f
C99 VOUT_SBCM VSS 1.66471f
C100 VOUT_RCCM VSS 3.08137f
C101 VAUX VSS 16.1107f
C102 VIN VSS 2.05138f
C103 EN VSS 1.41253f
C104 VDD VSS 0.23404p
C105 a_6883_483# VSS 2.90137f
C106 a_6293_483# VSS 6.39712f
C107 a_5657_4411# VSS 8.54632f
C108 a_5777_8307# VSS 7.65736f
C109 a_1385_n5930# VSS 12.1715f
C110 a_595_n5930# VSS 4.51891f
C111 a_n195_n5930# VSS 7.79334f
C112 a_865_n5930# VSS 0.15972f
C113 a_75_n5930# VSS 0.03433f
C114 a_n715_n5930# VSS 0.03454f
C115 a_n1505_n5930# VSS 2.68739f
C116 a_n30270_3049# VSS 2.76443f
C117 a_n36440_3049# VSS 40.2369f
C118 a_n31010_3002# VSS 0.2556f
C119 a_n18208_5979# VSS 0.40915f
C120 a_n29950_3049# VSS 5.40042f
C121 a_n18728_5979# VSS 0.29335f
C122 a_n39492_5979# VSS 12.9545f
C123 a_n48062_5772# VSS 2.75305f
C124 a_n40012_5979# VSS 0.28827f
C125 a_n26898_5979# VSS 3.15784f
C126 a_n26898_12584# VSS 0.17393f
C127 a_n48182_5979# VSS 3.23215f
C128 a_n48182_12584# VSS 0.19383f
C129 a_n48062_12376# VSS 6.28119f
C130 w_n49368_5436# VSS 0.49536p
.ends

