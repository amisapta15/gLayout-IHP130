* NGSPICE file created from INPUT_STAGE.ext - technology: gf180mcuD

.subckt INPUT_STAGE VIN VDD VOUT_VIN VOUT_CCM VOUT_BCM VOUT_VCM EN
X0 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0.1236n ps=0.44472m w=10u l=2u
X1 VOUT_VCM VIN a_n1110_n1500# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X2 a_n1900_n1500# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X3 VOUT_VIN VIN a_1260_n1500# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X4 a_n320_n1500# a_n1900_n1500# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X5 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X6 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X7 a_n1900_n1500# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X8 VOUT_BCM VIN a_n320_n1500# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X9 a_n1900_n1500# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X10 VIN VIN a_n1900_n1500# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X11 a_n1110_n1500# a_n1900_n1500# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X12 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X13 a_470_n1500# a_n1900_n1500# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X14 a_n1900_n1500# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X15 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X16 VOUT_CCM VIN a_470_n1500# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X17 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X18 a_n1900_n1500# a_n1900_n1500# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X19 a_1260_n1500# a_n1900_n1500# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
C0 VOUT_VIN a_n1110_n1500# 0.13684f
C1 a_1260_n1500# a_n1110_n1500# 0.30103f
C2 VOUT_BCM VOUT_CCM 0.33028f
C3 VIN VOUT_VCM 0.63416f
C4 a_n1900_n1500# a_n1110_n1500# 1.80913f
C5 a_n320_n1500# VIN 0.63243f
C6 a_1260_n1500# EN 0.28741f
C7 VOUT_VIN a_470_n1500# 0.13662f
C8 a_470_n1500# a_1260_n1500# 0.80509f
C9 VOUT_VIN VDD 2.21442f
C10 VDD a_1260_n1500# 6.35462f
C11 EN a_n1900_n1500# 2.15734f
C12 a_470_n1500# a_n1900_n1500# 1.46461f
C13 VDD a_n1900_n1500# 44.9171f
C14 VOUT_BCM a_n1110_n1500# 0.17152f
C15 VOUT_VIN VIN 0.54995f
C16 a_1260_n1500# VIN 0.62105f
C17 VOUT_CCM a_n1110_n1500# 0.17047f
C18 a_n320_n1500# VOUT_VCM 2.30103f
C19 VIN a_n1900_n1500# 3.41485f
C20 a_470_n1500# VOUT_BCM 2.29847f
C21 a_470_n1500# VOUT_CCM 2.39829f
C22 VDD VOUT_BCM 1.12778f
C23 VDD VOUT_CCM 1.1279f
C24 VOUT_VIN VOUT_VCM 0.08091f
C25 a_1260_n1500# VOUT_VCM 0.10003f
C26 VOUT_VIN a_n320_n1500# 0.13558f
C27 a_n320_n1500# a_1260_n1500# 0.30154f
C28 VOUT_BCM VIN 0.62309f
C29 VIN VOUT_CCM 0.62193f
C30 a_n1900_n1500# VOUT_VCM 0.13364f
C31 EN a_n1110_n1500# 0.00563f
C32 a_n320_n1500# a_n1900_n1500# 1.46427f
C33 a_470_n1500# a_n1110_n1500# 0.34178f
C34 VDD a_n1110_n1500# 7.43338f
C35 a_470_n1500# EN 0.00915f
C36 VOUT_VIN a_1260_n1500# 2.35844f
C37 VDD EN 11.072f
C38 VDD a_470_n1500# 7.51371f
C39 VOUT_BCM VOUT_VCM 0.3303f
C40 VIN a_n1110_n1500# 2.86501f
C41 VOUT_CCM VOUT_VCM 0.09982f
C42 a_n320_n1500# VOUT_BCM 2.40482f
C43 VOUT_VIN a_n1900_n1500# 0.96309f
C44 a_1260_n1500# a_n1900_n1500# 2.37681f
C45 a_n320_n1500# VOUT_CCM 0.17025f
C46 a_470_n1500# VIN 0.62333f
C47 VDD VIN 14.5258f
C48 VOUT_VIN VOUT_BCM 0.08038f
C49 a_1260_n1500# VOUT_BCM 0.10042f
C50 VOUT_VIN VOUT_CCM 0.31084f
C51 a_1260_n1500# VOUT_CCM 2.29591f
C52 VOUT_VCM a_n1110_n1500# 2.41261f
C53 a_n320_n1500# a_n1110_n1500# 0.84535f
C54 VOUT_BCM a_n1900_n1500# 0.13521f
C55 a_n1900_n1500# VOUT_CCM 0.13973f
C56 a_470_n1500# VOUT_VCM 0.10043f
C57 a_n320_n1500# EN 0.0069f
C58 a_n320_n1500# a_470_n1500# 0.84407f
C59 VDD VOUT_VCM 1.21291f
C60 VDD a_n320_n1500# 7.43186f
C61 VOUT_VIN VSUBS 0.38142f
C62 VOUT_CCM VSUBS 0.15405f
C63 VOUT_BCM VSUBS 0.15363f
C64 VOUT_VCM VSUBS 0.28097f
C65 VIN VSUBS 2.45016f
C66 EN VSUBS 1.80875f
C67 VDD VSUBS 0.30456p
C68 a_1260_n1500# VSUBS 0.15844f
C69 a_470_n1500# VSUBS 0.03326f
C70 a_n320_n1500# VSUBS 0.03284f
C71 a_n1110_n1500# VSUBS 0.03295f
C72 a_n1900_n1500# VSUBS 3.20944f
.ends

