** sch_path: /foss/designs/gLayout-mahowalders/blocks/composite/regulated_cascoded_cmirror/xschem/Chipathon2025_pads/xschem/io_secondary_3p3_DC_tb.sch
**.subckt io_secondary_3p3_DC_tb
V1 DVDD GND 3
V2 VDD GND 3
V3 DVSS GND 0
V4 VSS GND 0
V5 PAD GND PWL(0 -10 500n 10 1u -10)
XIO1 DVSS DVDD VSS VDD PAD asig gf180mcu_fd_io__asig_5p0_extracted
XIO2 VDD to_gate asig VSS io_secondary_3p3
**** begin user architecture code

.include /foss/designs/gLayout-mahowalders/blocks/composite/regulated_cascoded_cmirror/xschem/Chipathon2025_pads/xschem/gf180mcu_fd_io.spice
.include /foss/designs/gLayout-mahowalders/blocks/composite/regulated_cascoded_cmirror/xschem/Chipathon2025_pads/xschem/gf180mcu_fd_io__asig_5p0_extracted.spice


.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice diode_typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical




.control
tran 1n 1u
plot V(PAD)+12 V(ASIG)+6 V(to_gate)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  Chipathon2025_pads/xschem/symbols/io_secondary_3p3/io_secondary_3p3.sym # of pins=4
** sym_path: /foss/designs/gLayout-mahowalders/blocks/composite/regulated_cascoded_cmirror/xschem/Chipathon2025_pads/xschem/symbols/io_secondary_3p3/io_secondary_3p3.sym
** sch_path: /foss/designs/gLayout-mahowalders/blocks/composite/regulated_cascoded_cmirror/xschem/Chipathon2025_pads/xschem/symbols/io_secondary_3p3/io_secondary_3p3.sch
.subckt io_secondary_3p3 VDD to_gate ASIG3V3 VSS


*.iopin VSS
*.iopin VDD
*.iopin to_gate
*.iopin ASIG3V3
XR1 to_gate ASIG3V3 VDD ppolyf_u r_width=16e-6 r_length=4e-6 m=1
D2 VSS to_gate diode_nd2ps_03v3 area='10u * 10u ' pj='2*10u + 2*10u ' m=4
D1 to_gate VDD diode_pd2nw_03v3 area='10u * 10u ' pj='2*10u + 2*10u ' m=4
.ends

.GLOBAL GND
.end
