| units: 0.5 tech: gf180mcuD format: MIT
x a_n6357_n2535# a_n3305_371# a_n6357_n2535# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-3184 y=371 nfet_03v3
x a_n6357_n2535# a_n3305_371# a_n6357_n2535# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-824 y=371 nfet_03v3
x a_n15047_n2535# VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-14136 y=371 pfet_03v3
x VIN a_n15047_n2535# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-12556 y=-2534 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-5948 y=-2534 pfet_03v3
x a_n6357_n2535# a_n3305_371# a_n6357_n2535# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=2125 y=371 nfet_03v3
x a_n3305_371# VSS a_n3305_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-824 y=-2134 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=15335 y=371 pfet_03v3
x a_3185_371# a_14407_n2535# VOUT VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=14527 y=-2534 pfet_03v3
x a_n15047_n2535# VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-9396 y=371 pfet_03v3
x VSS VSS VSS VSS d=185600,3432 l=200 w=1600 x=-3792 y=-2134 nfet_03v3
x a_6237_n2535# VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=6357 y=371 pfet_03v3
x a_n15047_n2535# VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-7816 y=371 pfet_03v3
x a_n6357_n2535# a_2865_371# a_3185_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=2985 y=371 nfet_03v3
x a_n3305_371# VSS a_2865_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=2985 y=-2134 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=5549 y=4069 pfet_03v3
x a_6237_n2535# VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=8727 y=371 pfet_03v3
x a_3185_371# a_6237_n2535# a_3185_371# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=13467 y=-2534 pfet_03v3
x a_n15047_n2535# VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-11766 y=371 pfet_03v3
x a_n3305_371# VSS a_n3305_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=945 y=-2134 nfet_03v3
x a_6237_n2535# VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=12677 y=371 pfet_03v3
x a_3185_371# a_6237_n2535# a_3185_371# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=9517 y=-2534 pfet_03v3
x VIN a_n15047_n2535# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-10976 y=-2534 pfet_03v3
x a_n3305_371# VSS a_n3305_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-3184 y=-2134 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-15734 y=4069 pfet_03v3
x a_n6357_n2535# a_n3305_371# a_n6357_n2535# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=945 y=371 nfet_03v3
x a_n3305_371# VSS a_n3305_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=2125 y=-2134 nfet_03v3
x a_6237_n2535# VDD a_14407_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=14527 y=371 pfet_03v3
x a_n3305_371# VSS a_n3305_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-2004 y=-2134 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=7165 y=4069 pfet_03v3
x VIN a_n15047_n2535# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-14926 y=-2534 pfet_03v3
x a_n6357_n2535# a_n3305_371# a_n6357_n2535# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-1414 y=371 nfet_03v3
x a_n3305_371# VSS a_n3305_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-234 y=-2134 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=5549 y=371 pfet_03v3
x a_6237_n2535# VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=10307 y=371 pfet_03v3
x a_3185_371# a_6237_n2535# a_3185_371# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=7937 y=-2534 pfet_03v3
x a_3185_371# a_6237_n2535# a_3185_371# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=11887 y=-2534 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-14118 y=4069 pfet_03v3
x a_n15047_n2535# VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-13346 y=371 pfet_03v3
x VIN a_n15047_n2535# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-13346 y=-2534 pfet_03v3
x VIN a_n15047_n2535# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-7816 y=-2534 pfet_03v3
x VSS VSS VSS VSS d=185600,3432 l=200 w=1600 x=3593 y=371 nfet_03v3
x a_n3305_371# VSS a_n3305_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=355 y=-2134 nfet_03v3
x a_3185_371# a_6237_n2535# a_3185_371# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=6357 y=-2534 pfet_03v3
x a_n6357_n2535# a_n3305_371# a_n6357_n2535# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-234 y=371 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=15335 y=-2534 pfet_03v3
x VIN a_n6877_n2535# a_n6357_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-6756 y=-2534 pfet_03v3
x VSS VSS VSS VSS d=185600,3432 l=200 w=1600 x=-3792 y=371 nfet_03v3
x a_n6357_n2535# a_n3305_371# a_n6357_n2535# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-2004 y=371 nfet_03v3
x a_6237_n2535# VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=7937 y=371 pfet_03v3
x a_6237_n2535# VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=11887 y=371 pfet_03v3
x a_n15047_n2535# VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-10976 y=371 pfet_03v3
x a_n15047_n2535# VDD a_n6877_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-6756 y=371 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-15734 y=371 pfet_03v3
x VIN a_n15047_n2535# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-11766 y=-2534 pfet_03v3
x a_n3305_371# VSS a_n3305_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-2594 y=-2134 nfet_03v3
x EN VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-14926 y=4069 pfet_03v3
x a_n15047_n2535# VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-8606 y=371 pfet_03v3
x VIN a_n15047_n2535# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-10186 y=-2534 pfet_03v3
x a_n3305_371# VSS a_n3305_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=1535 y=-2134 nfet_03v3
x a_6237_n2535# VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=7147 y=371 pfet_03v3
x a_n15047_n2535# VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-10186 y=371 pfet_03v3
x a_n3305_371# VSS a_n3305_371# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-1414 y=-2134 nfet_03v3
x a_6237_n2535# VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=11097 y=371 pfet_03v3
x EN VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=6357 y=4069 pfet_03v3
x a_n6357_n2535# a_n3305_371# a_n6357_n2535# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-2594 y=371 nfet_03v3
x VSS VSS VSS VSS d=185600,3432 l=200 w=1600 x=3593 y=-2134 nfet_03v3
x a_6237_n2535# VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=9517 y=371 pfet_03v3
x a_6237_n2535# VDD a_6237_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=13467 y=371 pfet_03v3
x a_3185_371# a_6237_n2535# a_3185_371# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=8727 y=-2534 pfet_03v3
x a_3185_371# a_6237_n2535# a_3185_371# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=10307 y=-2534 pfet_03v3
x a_3185_371# a_6237_n2535# a_3185_371# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=12677 y=-2534 pfet_03v3
x a_n15047_n2535# VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-12556 y=371 pfet_03v3
x VIN a_n15047_n2535# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-14136 y=-2534 pfet_03v3
x VIN a_n15047_n2535# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-8606 y=-2534 pfet_03v3
x a_n6357_n2535# a_n3305_371# a_n6357_n2535# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=355 y=371 nfet_03v3
x a_n6357_n2535# a_n3305_371# a_n6357_n2535# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=1535 y=371 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-15734 y=-2534 pfet_03v3
x a_3185_371# a_6237_n2535# a_3185_371# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=11097 y=-2534 pfet_03v3
x a_n15047_n2535# VDD a_n15047_n2535# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-14926 y=371 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-5948 y=371 pfet_03v3
x VIN a_n15047_n2535# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-9396 y=-2534 pfet_03v3
x a_3185_371# a_6237_n2535# a_3185_371# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=7147 y=-2534 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=5549 y=-2534 pfet_03v3
C a_n6357_n2535# a_n3305_371# 36.6
C VDD a_n6877_n2535# 3.1
C EN a_n6877_n2535# 0.0
C VOUT a_14407_n2535# 0.9
C a_n15047_n2535# VDD 48.7
C EN a_n15047_n2535# 0.7
C a_14407_n2535# VDD 3.1
C a_n6357_n2535# VIN 0.5
C a_3185_371# a_14407_n2535# 1.0
C a_3185_371# a_2865_371# 1.1
C VOUT VDD 1.5
C a_n6357_n2535# a_n6877_n2535# 0.9
C EN VDD 5.8
C VIN a_n6877_n2535# 1.0
C a_3185_371# VOUT 0.5
C a_n3305_371# a_2865_371# 0.5
C a_14407_n2535# a_6237_n2535# 1.0
C a_3185_371# VDD 15.5
C a_3185_371# EN 0.0
C a_n6357_n2535# a_n15047_n2535# 0.1
C VIN a_n15047_n2535# 29.5
C a_n6357_n2535# a_2865_371# 0.9
C VOUT a_6237_n2535# 0.1
C a_6237_n2535# VDD 48.7
C EN a_6237_n2535# 0.7
C a_n15047_n2535# a_n6877_n2535# 1.0
C a_3185_371# a_6237_n2535# 29.5
C a_n6357_n2535# VDD 1.8
C EN a_n6357_n2535# 0.0
C VIN VDD 15.2
C a_3185_371# a_n6357_n2535# 0.3
C VOUT0 0.4
R VOUT 123
C VIN0 2.7
R VIN 1998
C EN0 5.8
R EN 120
C VDD0 538.9
R VDD 26835
R VSS 4899
C a_14407_n2535#0 0.3
R a_14407_n2535# 260
C a_3185_371#0 4.9
R a_3185_371# 2090
C a_2865_371#0 2.8
R a_2865_371# 191
C a_n3305_371#0 40.2
R a_n3305_371# 2962
C a_n6357_n2535#0 12.9
R a_n6357_n2535# 2054
C a_n6877_n2535#0 0.2
R a_n6877_n2535# 260
C a_6237_n2535#0 3.3
R a_6237_n2535# 3505
C a_n15047_n2535#0 3.2
R a_n15047_n2535# 3505
