magic
tech gf180mcuD
magscale 1 10
timestamp 1757961865
<< nwell >>
rect -4500 -1176 4500 1176
<< pwell >>
rect -4676 1176 4676 1352
rect -4676 -1176 -4500 1176
rect 4500 -1176 4676 1176
rect -4676 -1352 4676 -1176
<< mvpsubdiff >>
rect -4644 1248 4644 1320
rect -4644 1204 -4572 1248
rect -4644 -1204 -4631 1204
rect -4585 -1204 -4572 1204
rect 4572 1204 4644 1248
rect -4644 -1248 -4572 -1204
rect 4572 -1204 4585 1204
rect 4631 -1204 4644 1204
rect 4572 -1248 4644 -1204
rect -4644 -1320 4644 -1248
<< mvnsubdiff >>
rect -4468 1131 4468 1144
rect -4468 1085 -4352 1131
rect -2296 1085 -2136 1131
rect -80 1085 80 1131
rect 2136 1085 2296 1131
rect 4352 1085 4468 1131
rect -4468 1072 4468 1085
rect -4468 1028 -4396 1072
rect -4468 -1028 -4455 1028
rect -4409 -1028 -4396 1028
rect -2252 1028 -2180 1072
rect -4468 -1072 -4396 -1028
rect -2252 -1028 -2239 1028
rect -2193 -1028 -2180 1028
rect -36 1028 36 1072
rect -2252 -1072 -2180 -1028
rect -36 -1028 -23 1028
rect 23 -1028 36 1028
rect 2180 1028 2252 1072
rect -36 -1072 36 -1028
rect 2180 -1028 2193 1028
rect 2239 -1028 2252 1028
rect 4396 1028 4468 1072
rect 2180 -1072 2252 -1028
rect 4396 -1028 4409 1028
rect 4455 -1028 4468 1028
rect 4396 -1072 4468 -1028
rect -4468 -1085 4468 -1072
rect -4468 -1131 -4352 -1085
rect -2296 -1131 -2136 -1085
rect -80 -1131 80 -1085
rect 2136 -1131 2296 -1085
rect 4352 -1131 4468 -1085
rect -4468 -1144 4468 -1131
<< mvpsubdiffcont >>
rect -4631 -1204 -4585 1204
rect 4585 -1204 4631 1204
<< mvnsubdiffcont >>
rect -4352 1085 -2296 1131
rect -2136 1085 -80 1131
rect 80 1085 2136 1131
rect 2296 1085 4352 1131
rect -4455 -1028 -4409 1028
rect -2239 -1028 -2193 1028
rect -23 -1028 23 1028
rect 2193 -1028 2239 1028
rect 4409 -1028 4455 1028
rect -4352 -1131 -2296 -1085
rect -2136 -1131 -80 -1085
rect 80 -1131 2136 -1085
rect 2296 -1131 4352 -1085
<< mvpdiode >>
rect -4324 987 -2324 1000
rect -4324 -987 -4311 987
rect -2337 -987 -2324 987
rect -4324 -1000 -2324 -987
rect -2108 987 -108 1000
rect -2108 -987 -2095 987
rect -121 -987 -108 987
rect -2108 -1000 -108 -987
rect 108 987 2108 1000
rect 108 -987 121 987
rect 2095 -987 2108 987
rect 108 -1000 2108 -987
rect 2324 987 4324 1000
rect 2324 -987 2337 987
rect 4311 -987 4324 987
rect 2324 -1000 4324 -987
<< mvpdiodec >>
rect -4311 -987 -2337 987
rect -2095 -987 -121 987
rect 121 -987 2095 987
rect 2337 -987 4311 987
<< metal1 >>
rect -4631 1261 4631 1307
rect -4631 1204 -4585 1261
rect 4585 1204 4631 1261
rect -4455 1085 -4352 1131
rect -2296 1085 -2136 1131
rect -80 1085 80 1131
rect 2136 1085 2296 1131
rect 4352 1085 4455 1131
rect -4455 1028 -4409 1085
rect -2239 1028 -2193 1085
rect -4322 -987 -4311 987
rect -2337 -987 -2326 987
rect -4455 -1085 -4409 -1028
rect -23 1028 23 1085
rect -2106 -987 -2095 987
rect -121 -987 -110 987
rect -2239 -1085 -2193 -1028
rect 2193 1028 2239 1085
rect 110 -987 121 987
rect 2095 -987 2106 987
rect -23 -1085 23 -1028
rect 4409 1028 4455 1085
rect 2326 -987 2337 987
rect 4311 -987 4322 987
rect 2193 -1085 2239 -1028
rect 4409 -1085 4455 -1028
rect -4455 -1131 -4352 -1085
rect -2296 -1131 -2136 -1085
rect -80 -1131 80 -1085
rect 2136 -1131 2296 -1085
rect 4352 -1131 4455 -1085
rect -4631 -1261 -4585 -1204
rect 4585 -1261 4631 -1204
rect -4631 -1307 4631 -1261
<< properties >>
string diode_pd2nw_06v0_5DG9HC parameters
string FIXED_BBOX 2216 -1108 4432 1108
string gencell diode_pd2nw_06v0
string library gf180mcu
string parameters w 10 l 10 area 100.0 peri 40.0 nx 4 ny 1 dummy 0 lmin 0.45 wmin 0.45 class diode elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 0 gbc 0 doverlap 1 full_metal 1 compatible {diode_pd2nw_03v3 diode_pd2nw_06v0}
<< end >>
