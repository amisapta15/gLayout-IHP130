* NGSPICE file created from INPUT_STAGE.ext - technology: gf180mcuD

.subckt INPUT_STAGE VIN VDD VOUT_CCM VOUT_BCM VOUT_VCM EN
X0 a_n1505_n1396# a_n1505_n1396# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X1 a_n1505_n1396# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X2 VIN VIN a_n1505_n1396# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X3 VOUT_CCM VIN a_865_n1396# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X4 a_75_n1396# a_n1505_n1396# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X5 a_n1505_n1396# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X6 a_n1505_n1396# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X7 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0.1116n ps=0.40232m w=10u l=2u
X8 a_n715_n1396# a_n1505_n1396# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X9 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X10 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X11 VOUT_VCM VIN a_n715_n1396# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X12 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X13 VOUT_BCM VIN a_75_n1396# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X14 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X15 a_865_n1396# a_n1505_n1396# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X16 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
C0 a_n715_n1396# EN 0.00664f
C1 VOUT_VCM a_75_n1396# 2.03168f
C2 a_75_n1396# a_865_n1396# 0.74423f
C3 a_n1505_n1396# VDD 31.4897f
C4 a_n715_n1396# VIN 2.59448f
C5 a_n1505_n1396# a_75_n1396# 1.38044f
C6 VOUT_BCM VOUT_CCM 0.31085f
C7 EN a_865_n1396# 0.21853f
C8 VIN VOUT_VCM 0.63325f
C9 VIN a_865_n1396# 0.62292f
C10 a_n715_n1396# VOUT_VCM 2.02854f
C11 EN a_n1505_n1396# 1.62501f
C12 a_n715_n1396# a_865_n1396# 0.30282f
C13 VOUT_CCM VDD 1.99803f
C14 VIN a_n1505_n1396# 2.98274f
C15 VOUT_CCM a_75_n1396# 0.13665f
C16 a_n715_n1396# a_n1505_n1396# 1.68766f
C17 VOUT_BCM VDD 0.97996f
C18 VOUT_VCM a_865_n1396# 0.10043f
C19 VOUT_BCM a_75_n1396# 2.02098f
C20 a_n1505_n1396# VOUT_VCM 0.13478f
C21 a_n1505_n1396# a_865_n1396# 2.19448f
C22 VIN VOUT_CCM 0.55089f
C23 a_75_n1396# VDD 6.35872f
C24 a_n715_n1396# VOUT_CCM 0.13688f
C25 VOUT_BCM VIN 0.62256f
C26 VOUT_BCM a_n715_n1396# 0.17152f
C27 EN VDD 7.30305f
C28 VOUT_VCM VOUT_CCM 0.08093f
C29 VOUT_CCM a_865_n1396# 1.98101f
C30 VIN VDD 10.2566f
C31 EN a_75_n1396# 0.00866f
C32 a_n715_n1396# VDD 6.34675f
C33 VIN a_75_n1396# 0.6318f
C34 a_n1505_n1396# VOUT_CCM 0.7907f
C35 a_n715_n1396# a_75_n1396# 0.78447f
C36 VOUT_BCM VOUT_VCM 0.3303f
C37 VOUT_BCM a_865_n1396# 2.02912f
C38 VOUT_BCM a_n1505_n1396# 0.13836f
C39 VOUT_VCM VDD 1.06408f
C40 a_865_n1396# VDD 5.40929f
C41 VOUT_CCM VSUBS 0.38142f
C42 VOUT_BCM VSUBS 0.15342f
C43 VOUT_VCM VSUBS 0.28097f
C44 VIN VSUBS 2.05138f
C45 EN VSUBS 1.41253f
C46 VDD VSUBS 0.23405p
C47 a_865_n1396# VSUBS 0.15972f
C48 a_75_n1396# VSUBS 0.03433f
C49 a_n715_n1396# VSUBS 0.03454f
C50 a_n1505_n1396# VSUBS 2.73114f
.ends

