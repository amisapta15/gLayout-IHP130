| units: 0.5 tech: gf180mcuD format: MIT
x a_n1505_n1396# VDD a_n1505_n1396# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1384 y=3300 pfet_03v3
x EN VDD a_n1505_n1396# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-199 y=8101 pfet_03v3
x VIN a_n1505_n1396# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1384 y=-1395 pfet_03v3
x VIN a_865_n1396# VOUT_CCM VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=985 y=-1395 pfet_03v3
x a_n1505_n1396# VDD a_75_n1396# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=195 y=3300 pfet_03v3
x EN VDD a_n1505_n1396# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-989 y=8101 pfet_03v3
x EN VDD a_n1505_n1396# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=590 y=8101 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1398 y=8101 pfet_03v3
x a_n1505_n1396# VDD a_n715_n1396# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-594 y=3300 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2192 y=3300 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2192 y=-1395 pfet_03v3
x VIN a_n715_n1396# VOUT_VCM VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-594 y=-1395 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1793 y=-1395 pfet_03v3
x VIN a_75_n1396# VOUT_BCM VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=195 y=-1395 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-1797 y=8101 pfet_03v3
x a_n1505_n1396# VDD a_865_n1396# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=985 y=3300 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1793 y=3300 pfet_03v3
C VIN VDD 10.3
C VOUT_BCM a_n715_n1396# 0.2
C a_n1505_n1396# VOUT_VCM 0.1
C a_865_n1396# a_n715_n1396# 0.3
C VOUT_BCM VDD 1.0
C a_n715_n1396# a_75_n1396# 0.8
C a_n1505_n1396# EN 1.6
C VOUT_CCM VIN 0.6
C a_865_n1396# VDD 5.4
C a_n715_n1396# VOUT_VCM 2.0
C a_75_n1396# VDD 6.4
C VOUT_BCM VOUT_CCM 0.3
C VDD VOUT_VCM 1.1
C a_865_n1396# VOUT_CCM 2.0
C VOUT_BCM VIN 0.6
C a_n715_n1396# EN 0.0
C VOUT_CCM a_75_n1396# 0.1
C a_n1505_n1396# a_n715_n1396# 1.7
C a_865_n1396# VIN 0.6
C VDD EN 7.3
C VOUT_CCM VOUT_VCM 0.1
C a_n1505_n1396# VDD 31.5
C a_75_n1396# VIN 0.6
C a_865_n1396# VOUT_BCM 2.0
C VIN VOUT_VCM 0.6
C VOUT_BCM a_75_n1396# 2.0
C a_n1505_n1396# VOUT_CCM 0.8
C a_865_n1396# a_75_n1396# 0.7
C VOUT_BCM VOUT_VCM 0.3
C a_n715_n1396# VDD 6.3
C a_865_n1396# VOUT_VCM 0.1
C a_n1505_n1396# VIN 3.0
C a_75_n1396# VOUT_VCM 2.0
C VOUT_BCM a_n1505_n1396# 0.1
C VOUT_CCM a_n715_n1396# 0.1
C a_865_n1396# EN 0.2
C a_865_n1396# a_n1505_n1396# 2.2
C VOUT_CCM VDD 2.0
C a_75_n1396# EN 0.0
C a_n715_n1396# VIN 2.6
C a_n1505_n1396# a_75_n1396# 1.4
C VOUT_CCM0 0.4
R VOUT_CCM 127
C VOUT_BCM0 0.2
R VOUT_BCM 127
C VOUT_VCM0 0.3
R VOUT_VCM 127
C VIN0 2.1
R VIN 414
C EN0 1.4
R EN 198
C VDD0 234.1
R VDD 9009
C a_865_n1396#0 0.2
R a_865_n1396# 269
C a_75_n1396#0 0.0
R a_75_n1396# 269
C a_n715_n1396#0 0.0
R a_n715_n1396# 269
C a_n1505_n1396#0 2.7
R a_n1505_n1396# 974
