** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/buffer_tb.sch
**.subckt buffer_tb
Vdd net1 GND 1.65
Vin in GND dc 0 ac 0 pulse(0, 1.65, 0, 100p, 100p, 2n, 4n )
xinv1 net1 in out GND inv
xbuff1 net1 out outB GND buff
* noconn outB
**** begin user architecture code


.param temp=27

.control
save all
tran 50p 20n

* plot waveforms
plot v(in) v(out) v(outB)
.endc



 .lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ_stat

**** end user architecture code
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/inv.sym
** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/inv.sch
.subckt inv VDD in out VSS
*.iopin VDD
*.ipin in
*.iopin VSS
*.opin out
XM1 out in VSS VSS sg13_lv_nmos w=2.0u l=0.28u ng=1 m=1
XM2 out in VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=1
.ends


* expanding   symbol:  buff.sym # of pins=4
** sym_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/buff.sym
** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/buff.sch
.subckt buff VDD in out VSS
*.iopin VDD
*.ipin in
*.iopin VSS
*.opin out
XM1 net1 in VSS VSS sg13_lv_nmos w=0.5u l=0.28u ng=1 m=1
XM2 net1 in VDD VDD sg13_lv_pmos w=0.5u l=0.28u ng=2 m=1
XM4 out net1 VSS VSS sg13_lv_nmos w=0.87u l=0.28u ng=4 m=1
XM5 out net1 VDD VDD sg13_lv_pmos w=1.5u l=0.28u ng=4 m=1
.ends

.GLOBAL GND
.end
