* Extracted by KLayout with GF180MCU LVS runset on : 26/09/2025 14:50

.SUBCKT TOP VSS VDD PD|Z|tieH EN PU|ZN|tieL VBIAS VCM_OUT VIN_OUT BCM_OUT
+ CCM_OUT VIN gf180mcu_gnd
M$1 VDD VDD VDD VDD pfet_03v3 L=2U W=180U AS=104.4P AD=104.4P PS=380.88U
+ PD=380.88U
M$2 \$317 \$317 \$265 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$3 \$248 \$317 \$247 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$4 \$250 \$317 \$249 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$5 \$252 \$317 \$251 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$6 VIN_OUT \$317 \$253 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$9 \$265 \$265 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$10 \$247 \$265 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$11 \$249 \$265 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$12 \$251 \$265 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$13 \$253 \$265 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$16 \$222 \$222 \$354 VDD pfet_03v3 L=2U W=100U AS=60P AD=60P PS=212U PD=212U
M$26 \$356 \$222 \$355 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$29 \$347 \$347 \$358 VDD pfet_03v3 L=2U W=100U AS=60P AD=60P PS=212U PD=212U
M$39 \$314 \$347 \$359 VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$42 \$265 \$149 VDD VDD pfet_03v3 L=2U W=40U AS=24P AD=24P PS=84.8U PD=84.8U
M$48 \$354 \$354 VDD VDD pfet_03v3 L=2U W=100U AS=60P AD=60P PS=212U PD=212U
M$58 \$355 \$354 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$61 \$358 \$358 VDD VDD pfet_03v3 L=2U W=100U AS=60P AD=60P PS=212U PD=212U
M$71 \$359 \$358 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$74 \$354 \$149 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$77 \$358 \$149 VDD VDD pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U PD=21.2U
M$79 \$202 \$202 VDD VDD pfet_05v0 L=0.5U W=0.9U AS=0.396P AD=0.396P PS=2.68U
+ PD=2.68U
M$80 PD|Z|tieH \$207 VDD VDD pfet_05v0 L=0.5U W=0.9U AS=0.396P AD=0.396P
+ PS=2.68U PD=2.68U
M$81 VSS VSS VSS gf180mcu_gnd nfet_03v3 L=1U W=32U AS=18.56P AD=18.56P
+ PS=68.64U PD=68.64U
M$82 \$357 \$357 VSS gf180mcu_gnd nfet_03v3 L=1U W=80U AS=48P AD=48P PS=172U
+ PD=172U
M$92 \$368 \$357 VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P PS=17.2U
+ PD=17.2U
M$95 \$356 \$356 \$357 gf180mcu_gnd nfet_03v3 L=1U W=80U AS=48P AD=48P PS=172U
+ PD=172U
M$105 \$347 \$356 \$368 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$107 PU|ZN|tieL \$202 VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.66U AS=0.2904P
+ AD=0.2904P PS=2.2U PD=2.2U
M$108 \$207 \$207 VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.66U AS=0.2904P
+ AD=0.2904P PS=2.2U PD=2.2U
M$109 VSS VSS VSS VSS nfet_03v3_dn L=1U W=48U AS=27.84P AD=27.84P PS=109.92U
+ PD=109.92U
M$110 \$248 \$248 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$111 VCM_OUT \$248 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$114 \$268 \$268 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$115 \$288 \$268 VSS VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U PD=9.2U
M$118 \$250 \$250 \$268 VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$119 BCM_OUT \$250 \$288 VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$122 CCM_OUT \$314 \$312 VSS nfet_03v3_dn L=1U W=8U AS=4.8P AD=4.8P PS=18.4U
+ PD=18.4U
M$123 \$314 \$312 VSS VSS nfet_03v3_dn L=1U W=8U AS=4.8P AD=4.8P PS=18.4U
+ PD=18.4U
M$128 \$348 \$252 VSS VSS nfet_03v3_dn L=1U W=8U AS=4.8P AD=4.8P PS=18.4U
+ PD=18.4U
M$129 \$312 \$252 VSS VSS nfet_03v3_dn L=1U W=8U AS=4.8P AD=4.8P PS=18.4U
+ PD=18.4U
M$134 \$314 \$348 VSS VSS nfet_03v3_dn L=1U W=8U AS=4.8P AD=4.8P PS=18.4U
+ PD=18.4U
M$135 \$252 \$314 \$348 VSS nfet_03v3_dn L=1U W=8U AS=4.8P AD=4.8P PS=18.4U
+ PD=18.4U
D$139 VSS \$149 diode_nd2ps_06v0 A=400P P=160U
D$143 VSS \$222 diode_nd2ps_06v0 A=400P P=160U
D$147 VSS \$317 diode_nd2ps_06v0 A=400P P=160U
D$151 \$149 VDD diode_pd2nw_06v0 A=400P P=160U
D$155 \$222 VDD diode_pd2nw_06v0 A=400P P=160U
D$159 \$317 VDD diode_pd2nw_06v0 A=400P P=160U
R$163 \$149 EN gf180mcu_gnd 87.5 ppolyf_u L=10U W=40U
R$164 \$222 VBIAS gf180mcu_gnd 87.5 ppolyf_u L=10U W=40U
R$165 \$317 VIN gf180mcu_gnd 87.5 ppolyf_u L=10U W=40U
.ENDS TOP
