* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VIN VSS VDD VOUT_RCCM VOUT_SBCM VOUT_VCM VAUX EN
X0 VAUX a_5777_8307# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X1 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X2 VAUX a_5777_8307# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X3 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0.17441n ps=0.65676m w=4u l=1u
X4 VAUX a_5657_4411# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X5 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X6 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X7 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X8 a_n40012_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X9 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X10 VAUX a_5657_4411# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X11 a_n715_n5930# a_n1505_n5930# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X12 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0.1116n ps=0.40232m w=10u l=2u
X13 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X14 a_n30270_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X15 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X16 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X17 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X18 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X19 a_n195_n5930# VIN a_n715_n5930# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X20 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X21 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X22 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X23 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X24 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X25 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X26 a_75_n5930# a_n1505_n5930# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X27 a_595_n5930# a_595_n5930# a_6293_483# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X28 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X29 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X30 a_1385_n5930# VAUX a_5777_8307# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X31 a_1385_n5930# VAUX a_5777_8307# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X32 a_595_n5930# VIN a_75_n5930# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X33 a_n1505_n5930# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X34 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X35 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X36 a_n29950_3049# a_n39492_5979# a_n30270_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X37 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X38 a_6883_483# a_6293_483# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X39 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X40 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0.27118n ps=0.97416m w=10u l=2u
X41 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X42 a_5777_8307# a_1385_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X43 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X44 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X45 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X46 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X47 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.7971p pd=21.15u as=0 ps=0 w=9.995u l=2u
X48 a_5777_8307# a_1385_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X49 a_n18208_5979# a_n29950_3049# a_n18728_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X50 VOUT_VCM a_n195_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X51 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X52 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X53 VOUT_SBCM a_595_n5930# a_6883_483# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X54 VSS VSS VSS VSS nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X55 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X56 a_n26898_5979# a_n48062_12376# a_n26898_12584# w_n49368_5436# pfet_03v3 ad=5.997p pd=21.19u as=5.997p ps=21.19u w=9.995u l=2u
X57 VSS VSS VSS VSS nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X58 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X59 a_n48182_5979# a_n48062_12376# a_n48182_12584# w_n49368_5436# pfet_03v3 ad=5.997p pd=21.19u as=5.997p ps=21.19u w=9.995u l=2u
X60 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X61 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X62 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X63 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X64 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X65 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X66 a_5657_4411# a_1385_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X67 a_5657_4411# a_1385_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X68 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X69 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X70 VSS VSS VSS VSS nfet_03v3 ad=4.6429p pd=17.17u as=0 ps=0 w=8.005u l=1u
X71 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X72 a_n39492_5979# a_n48062_5772# a_n40012_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X73 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X74 a_n1505_n5930# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X75 a_n1505_n5930# a_n1505_n5930# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X76 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X77 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X78 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X79 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X80 a_n39492_5979# a_n31010_3002# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X81 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X82 VIN VIN a_n1505_n5930# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X83 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X84 a_n1505_n5930# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X85 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X86 a_865_n5930# a_n1505_n5930# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X87 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X88 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X89 a_6293_483# a_6293_483# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X90 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X91 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X92 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X93 a_1385_n5930# VIN a_865_n5930# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X94 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X95 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X96 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X97 a_n195_n5930# a_n195_n5930# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X98 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X99 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X100 a_n29950_3049# a_n29950_3049# a_n26898_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X101 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X102 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X103 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X104 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X105 a_n18728_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X106 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.7971p pd=21.15u as=0 ps=0 w=9.995u l=2u
X107 VOUT_RCCM VAUX a_5657_4411# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X108 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X109 VSS VSS VSS VSS nfet_03v3 ad=4.6429p pd=17.17u as=0 ps=0 w=8.005u l=1u
X110 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X111 VOUT_RCCM VAUX a_5657_4411# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X112 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X113 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.7971p pd=21.15u as=0 ps=0 w=9.995u l=2u
X114 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X115 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.7971p pd=21.15u as=0 ps=0 w=9.995u l=2u
X116 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X117 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X118 a_n36440_3049# a_n36440_3049# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X119 a_n39492_5979# a_n39492_5979# a_n36440_3049# VSS nfet_03v3 ad=4.803p pd=17.21u as=4.803p ps=17.21u w=8.005u l=1u
X120 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X121 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X122 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X123 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X124 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X125 a_n48062_5772# a_n48062_5772# a_n48182_5979# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X126 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X127 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X128 a_n48182_5979# a_n48182_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X129 a_n26898_5979# a_n26898_5979# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X130 w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
.ends

