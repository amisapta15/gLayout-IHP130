* NGSPICE file created from RCM.ext - technology: gf180mcuD

.subckt RCM VIN VSS VAUX VOUT
X0 VAUX a_n985_3311# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X1 a_n1105_n585# VIN VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X2 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=47.04p ps=0.18352m w=4u l=1u
X3 a_n985_3311# VIN VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X4 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X5 VOUT VAUX a_n1105_n585# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X6 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X7 VAUX a_n985_3311# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X8 VAUX a_n1105_n585# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X9 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X10 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X11 VIN VAUX a_n985_3311# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X12 VAUX a_n1105_n585# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X13 a_n985_3311# VIN VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X14 VIN VAUX a_n985_3311# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X15 VOUT VAUX a_n1105_n585# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X16 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X17 a_n1105_n585# VIN VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
C0 VAUX a_n985_3311# 3.58908f
C1 a_n985_3311# a_n1105_n585# 0.36393f
C2 VIN a_n985_3311# 3.00275f
C3 VOUT a_n985_3311# 0.0136f
C4 VAUX a_n1105_n585# 3.29507f
C5 VAUX VIN 1.44115f
C6 VOUT VAUX 0.57679f
C7 VIN a_n1105_n585# 0.85546f
C8 VOUT a_n1105_n585# 2.17202f
C9 VOUT VIN 0.00933f
C10 VOUT VSS 3.08137f
C11 VIN VSS 7.81372f
C12 VAUX VSS 12.7612f
C13 a_n1105_n585# VSS 8.53412f
C14 a_n985_3311# VSS 7.65736f
.ends

