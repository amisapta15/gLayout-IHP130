| units: 0.5 tech: gf180mcuD format: MIT
x a_n985_3311# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=195 y=3691 nfet_03v3
x VIN VSS a_n1105_n585# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=785 y=1553 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=-1592 y=-584 nfet_03v3
x VIN VSS a_n985_3311# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=195 y=1553 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=-1592 y=3691 nfet_03v3
x VAUX a_n1105_n585# VOUT VSS s=96000,1840 d=96000,1840 l=200 w=800 x=-984 y=-584 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=1393 y=-584 nfet_03v3
x a_n985_3311# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=-984 y=3691 nfet_03v3
x a_n1105_n585# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=-394 y=-584 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=1393 y=3691 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=-1592 y=1553 nfet_03v3
x VAUX a_n985_3311# VIN VSS s=96000,1840 d=96000,1840 l=200 w=800 x=-394 y=3691 nfet_03v3
x a_n1105_n585# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=785 y=-584 nfet_03v3
x VIN VSS a_n985_3311# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=-984 y=1553 nfet_03v3
x VAUX a_n985_3311# VIN VSS s=96000,1840 d=96000,1840 l=200 w=800 x=785 y=3691 nfet_03v3
x VAUX a_n1105_n585# VOUT VSS s=96000,1840 d=96000,1840 l=200 w=800 x=195 y=-584 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=1393 y=1553 nfet_03v3
x VIN VSS a_n1105_n585# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=-394 y=1553 nfet_03v3
C VAUX a_n985_3311# 3.6
C VAUX a_n1105_n585# 3.3
C VAUX VOUT 0.6
C VAUX VIN 1.4
C a_n1105_n585# a_n985_3311# 0.4
C VOUT a_n985_3311# 0.0
C VIN a_n985_3311# 3.0
C a_n1105_n585# VOUT 2.2
C a_n1105_n585# VIN 0.9
C VIN VOUT 0.0
C VOUT0 3.1
R VOUT 107
C VIN0 7.8
R VIN 347
C VAUX0 12.8
R VAUX 469
R VSS 3589
C a_n1105_n585#0 8.5
R a_n1105_n585# 340
C a_n985_3311#0 7.7
R a_n985_3311# 335
