| units: 0.5 tech: gf180mcuD format: MIT
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=-1002 y=-584 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=803 y=-584 nfet_03v3
x VIN VSS VIN VSS s=96000,1840 d=96000,1840 l=200 w=800 x=-394 y=-584 nfet_03v3
x VIN VSS VOUT VSS s=96000,1840 d=96000,1840 l=200 w=800 x=195 y=-584 nfet_03v3
C VOUT VIN 0.2
C VOUT0 3.0
R VOUT 47
C VIN0 5.9
R VIN 159
R VSS 1473
