* NGSPICE file created from M.ext - technology: sky130A

.subckt M VIN VSS VDD VOUT_VIN VOUT_RCCM VOUT_SBCM VOUT_VCM VAUX EN
X0 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X1 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=115.44 ps=634.90002 w=4 l=1
X2 a_n17107_9910# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X3 a_200_n5640# a_200_n5640# a_6260_503# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X4 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X5 VOUT_RCCM a_5835_4440# a_5757_4829# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X6 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=81.9078 ps=436.42001 w=10 l=2
X7 a_n32245_7124# EN w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X8 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X9 a_6722_503# a_6260_503# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X10 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X11 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X12 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X13 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X14 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X15 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X16 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X17 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X18 a_5835_4440# a_5757_4829# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X19 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X20 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X21 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=0 ps=0 w=10.005 l=2
X22 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=187.2 ps=997.44 w=10 l=2
X23 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=0 ps=0 w=10.005 l=2
X24 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X25 a_n1602_n5640# EN w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X26 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X27 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X28 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X29 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X30 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X31 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X32 a_5835_8163# a_862_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X33 a_n1602_n5640# EN w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X34 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X35 VOUT_VCM a_n462_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X36 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X37 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X38 a_5757_4829# a_862_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X39 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X40 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X41 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X42 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X43 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X44 a_5835_4440# a_5835_8163# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X45 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X46 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X47 a_n278_n5640# a_n1602_n5640# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X48 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X49 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X50 a_1046_n5640# a_n1602_n5640# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X51 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X52 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X53 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X54 a_200_n5640# a_n1524_n6691# a_n278_n5640# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=3.90195 ps=20.79 w=10.005 l=2
X55 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X56 a_384_n5640# a_n1602_n5640# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X57 a_862_n5640# a_5835_4440# a_5835_8163# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X58 a_6260_503# a_6260_503# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X59 a_n6641_7124# a_n16829_9910# a_n7119_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X60 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X61 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X62 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X63 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X64 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X65 a_n1602_n5640# EN w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X66 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X67 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X68 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X69 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X70 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X71 VOUT_VIN a_n1524_n6691# a_1046_n5640# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=3.90195 ps=20.79 w=10.005 l=2
X72 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X73 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X74 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X75 a_n24817_7124# VAUX a_n25295_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X76 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X77 VOUT_RCCM a_5835_4440# a_5757_4829# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X78 a_n462_n5640# a_n462_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X79 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X80 a_5835_4440# a_5757_4829# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X81 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X82 a_n1524_n6691# a_n1524_n6691# a_n1602_n5640# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=3.90195 ps=20.79 w=10.005 l=2
X83 a_n940_n5640# a_n1602_n5640# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X84 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X85 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X86 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X87 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X88 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X89 a_n1602_n5640# a_n1602_n5640# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X90 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X91 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X92 a_n16829_9910# a_n24817_7124# a_n17107_9910# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X93 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X94 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X95 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X96 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X97 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X98 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X99 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X100 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X101 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X102 a_5835_8163# a_862_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X103 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X104 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X105 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X106 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X107 a_5757_4829# a_862_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X108 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X109 a_n7119_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X110 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X111 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X112 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X113 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X114 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X115 VOUT_SBCM a_200_n5640# a_6722_503# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X116 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X117 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X118 a_5835_4440# a_5835_8163# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X119 a_n462_n5640# a_n1524_n6691# a_n940_n5640# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=3.90195 ps=20.79 w=10.005 l=2
X120 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X121 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X122 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X123 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X124 a_n25295_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X125 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X126 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X127 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X128 a_862_n5640# a_5835_4440# a_5835_8163# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X129 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X130 a_862_n5640# a_n1524_n6691# a_384_n5640# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=3.90195 ps=20.79 w=10.005 l=2
X131 a_n14069_7124# EN w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X132 a_n1602_n5640# EN w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X133 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
C0 a_n22057_9909# a_n24817_7124# 36.2281f
C1 a_n940_n5640# a_n278_n5640# 0.67164f
C2 a_5835_8163# a_5757_4829# 0.30219f
C3 li_n5290_9325# a_862_n5640# 0.06369f
C4 li_n32467_15897# EN 0.00835f
C5 li_n3142_n10147# li_9474_n10147# 0.04039f
C6 EN li_n5290_9325# 0.04046f
C7 a_1046_n5640# a_384_n5640# 0.63691f
C8 a_384_n5640# a_862_n5640# 2.34599f
C9 VAUX w_n33347_6533# 15.0569f
C10 w_n2704_n7119# a_n1602_n5640# 43.9057f
C11 a_n22057_9909# a_n17107_9910# 0.66142f
C12 EN a_n32245_7124# 1.1821f
C13 a_200_n5640# a_n1602_n5640# 0.1065f
C14 a_5835_4440# a_5757_4829# 3.29564f
C15 EN a_384_n5640# 0.0053f
C16 a_6260_503# a_200_n5640# 1.83044f
C17 w_n2704_n7119# w_n33347_6533# 4.70379f
C18 a_n1524_n6691# a_n278_n5640# 0.87226f
C19 VOUT_VIN w_n2704_n7119# 2.58391f
C20 VOUT_VIN a_200_n5640# 0.06549f
C21 a_5835_8163# li_6128_10166# 0.00509f
C22 EN a_n7119_7124# 0
C23 a_5835_8163# a_862_n5640# 2.8133f
C24 a_n25295_7124# a_n32245_7124# 1.36306f
C25 a_1046_n5640# a_n1602_n5640# 2.67319f
C26 w_n2704_n7119# VAUX 0.04078f
C27 a_862_n5640# a_n1602_n5640# 0.42329f
C28 a_5835_4440# li_6128_10166# 0.00115f
C29 a_n462_n5640# a_384_n5640# 0.08474f
C30 li_9462_n10101# li_9474_n10147# 0.04039f
C31 li_9462_n10101# VOUT_VIN 0.06234f
C32 VOUT_VIN li_6128_10166# 0.7554f
C33 a_5835_4440# a_862_n5640# 1.45234f
C34 EN a_n1602_n5640# 3.24529f
C35 li_n32467_15897# VDD 0.05752f
C36 w_n2704_n7119# a_200_n5640# 0.98885f
C37 a_n7119_7124# a_n16829_9910# 1.17654f
C38 VOUT_VIN a_1046_n5640# 2.3704f
C39 VOUT_VIN a_862_n5640# 2.97221f
C40 EN w_n33347_6533# 6.7823f
C41 a_n940_n5640# a_384_n5640# 0.29693f
C42 VOUT_RCCM a_5835_8163# 0.00529f
C43 a_n16829_9910# a_n24817_7124# 0.48217f
C44 li_9462_n10101# VAUX 0.04046f
C45 a_n25295_7124# a_n24817_7124# 0.81434f
C46 VAUX li_6128_10166# 0.48902f
C47 VSS li_6128_10166# 0.08424f
C48 a_n17107_9910# a_n16829_9910# 0.94941f
C49 a_5835_4440# VOUT_RCCM 0.73487f
C50 a_862_n5640# a_5757_4829# 1.12178f
C51 a_n462_n5640# a_n1602_n5640# 0.10518f
C52 VAUX EN 0.00277f
C53 w_n2704_n7119# a_1046_n5640# 5.82159f
C54 a_n6641_7124# a_n16829_9910# 0.77125f
C55 a_200_n5640# a_1046_n5640# 0.08447f
C56 w_n2704_n7119# a_862_n5640# 1.65196f
C57 a_200_n5640# a_862_n5640# 0.34342f
C58 a_n16829_9910# w_n33347_6533# 14.6684f
C59 a_n1524_n6691# a_384_n5640# 0.86491f
C60 a_n25295_7124# w_n33347_6533# 2.9256f
C61 a_n278_n5640# a_384_n5640# 0.67118f
C62 w_n2704_n7119# EN 13.8092f
C63 VOUT_SBCM a_6722_503# 1.00834f
C64 VOUT_VIN a_n462_n5640# 0.06623f
C65 a_n14069_7124# a_n7119_7124# 1.36306f
C66 a_n940_n5640# a_n1602_n5640# 2.26345f
C67 VOUT_RCCM a_5757_4829# 1.83249f
C68 VOUT_VIN a_n940_n5640# 0.12116f
C69 VAUX a_n25295_7124# 1.17654f
C70 a_1046_n5640# a_862_n5640# 1.88942f
C71 li_9462_n10101# EN 0.06634f
C72 w_n2704_n7119# a_n16829_9910# 0.04377f
C73 EN li_6128_10166# 0.78481f
C74 w_n2704_n7119# a_n462_n5640# 1.08876f
C75 a_n1524_n6691# a_n1602_n5640# 3.76054f
C76 EN a_1046_n5640# 0.23129f
C77 a_n14069_7124# a_n6641_7124# 0.04849f
C78 a_200_n5640# a_n462_n5640# 0.65327f
C79 a_n278_n5640# a_n1602_n5640# 1.98713f
C80 a_n14069_7124# w_n33347_6533# 48.675f
C81 li_9462_n10101# VIN 0.041f
C82 li_n32467_15897# a_n32245_7124# 0.00846f
C83 li_9462_n10101# VOUT_RCCM 0.0631f
C84 VOUT_VIN a_n1524_n6691# 0.81264f
C85 a_n940_n5640# w_n2704_n7119# 6.63356f
C86 VOUT_VIN a_n278_n5640# 0.12086f
C87 a_n940_n5640# a_200_n5640# 0.14873f
C88 VOUT_RCCM a_862_n5640# 0.0044f
C89 li_n3142_n10147# a_n1524_n6691# 0.04745f
C90 a_n462_n5640# a_1046_n5640# 0.08404f
C91 a_n462_n5640# a_862_n5640# 0.08458f
C92 a_n7119_7124# li_n5290_9325# 0
C93 EN a_n25295_7124# 0
C94 w_n2704_n7119# a_n1524_n6691# 14.2578f
C95 VOUT_SBCM a_6260_503# 0.06811f
C96 a_6260_503# a_6722_503# 0.42557f
C97 a_n1524_n6691# a_200_n5640# 0.86559f
C98 w_n2704_n7119# a_n278_n5640# 6.62307f
C99 a_n278_n5640# a_200_n5640# 2.35168f
C100 a_n940_n5640# a_1046_n5640# 0.26163f
C101 a_n940_n5640# a_862_n5640# 0.14828f
C102 a_n24817_7124# a_n32245_7124# 0.05105f
C103 a_n940_n5640# EN 0.00394f
C104 li_n32467_15897# w_n33347_6533# 1.08918f
C105 li_n5290_9325# a_n6641_7124# 0.03696f
C106 a_5835_4440# li_n5290_9325# 0.04254f
C107 li_n5290_9325# w_n33347_6533# 0.02663f
C108 a_384_n5640# a_n1602_n5640# 1.98675f
C109 VOUT_VIN li_n5290_9325# 0.06228f
C110 a_n1524_n6691# a_1046_n5640# 0.86259f
C111 a_n32245_7124# w_n33347_6533# 48.687f
C112 a_n278_n5640# a_1046_n5640# 0.26233f
C113 a_n1524_n6691# a_862_n5640# 0.86245f
C114 a_n278_n5640# a_862_n5640# 0.14816f
C115 a_n14069_7124# EN 1.18736f
C116 VOUT_SBCM a_200_n5640# 0.29896f
C117 li_n32467_15897# VAUX 0.51079f
C118 a_6722_503# a_200_n5640# 1.27665f
C119 VOUT_VCM li_9462_n10101# 0.06295f
C120 VOUT_VIN a_384_n5640# 0.12131f
C121 a_n278_n5640# EN 0.00433f
C122 a_n940_n5640# a_n462_n5640# 2.37036f
C123 a_n7119_7124# a_n6641_7124# 0.75352f
C124 a_n7119_7124# w_n33347_6533# 2.9256f
C125 a_n17107_9910# a_n24817_7124# 1.04802f
C126 VAUX a_n32245_7124# 30.6991f
C127 a_n24817_7124# w_n33347_6533# 1.6542f
C128 a_5835_4440# a_5835_8163# 3.63338f
C129 a_n14069_7124# a_n16829_9910# 30.6918f
C130 li_9462_n10101# VOUT_SBCM 0.06295f
C131 VOUT_VIN a_5835_8163# 0
C132 w_n2704_n7119# a_384_n5640# 6.70512f
C133 a_200_n5640# a_384_n5640# 1.88756f
C134 a_n1524_n6691# a_n462_n5640# 0.87278f
C135 a_n278_n5640# a_n462_n5640# 1.89721f
C136 a_n17107_9910# w_n33347_6533# 0
C137 VOUT_VIN a_n1602_n5640# 0.62032f
C138 a_n6641_7124# w_n33347_6533# 1.39143f
C139 VAUX a_n24817_7124# 0.77125f
C140 VOUT_VIN a_5835_4440# 0.1026f
C141 VOUT_VCM a_n462_n5640# 0.30117f
C142 a_n940_n5640# a_n1524_n6691# 2.70328f
C143 VIN a_n22897_6995# 0.0814f
C144 VSS a_n22897_6995# 0.14776f
C145 VDD a_n22897_6995# 0.08953f
C146 VOUT_VCM a_n22897_6995# 5.45532f
C147 VOUT_VIN a_n22897_6995# 10.2333f
C148 VOUT_SBCM a_n22897_6995# 4.24238f
C149 VOUT_RCCM a_n22897_6995# 5.27364f
C150 VAUX a_n22897_6995# 25.2961f
C151 EN a_n22897_6995# 22.9185f
C152 li_9474_n10147# a_n22897_6995# 0.04374f $ **FLOATING
C153 li_n3142_n10147# a_n22897_6995# 5.84569f $ **FLOATING
C154 li_n5290_9325# a_n22897_6995# 4.6163f $ **FLOATING
C155 li_9462_n10101# a_n22897_6995# 18.8662f $ **FLOATING
C156 li_6128_10166# a_n22897_6995# 41.0831f $ **FLOATING
C157 li_n32467_15897# a_n22897_6995# 92.0531f $ **FLOATING
C158 a_n462_n5640# a_n22897_6995# 7.85547f
C159 a_n1524_n6691# a_n22897_6995# 4.10409f
C160 a_6722_503# a_n22897_6995# 2.58243f
C161 a_6260_503# a_n22897_6995# 6.07815f
C162 a_200_n5640# a_n22897_6995# 5.03421f
C163 a_1046_n5640# a_n22897_6995# 0.01985f
C164 a_5757_4829# a_n22897_6995# 7.57342f
C165 a_n1602_n5640# a_n22897_6995# 2.1896f
C166 a_862_n5640# a_n22897_6995# 11.9689f
C167 a_5835_4440# a_n22897_6995# 11.702f
C168 a_5835_8163# a_n22897_6995# 6.91168f
C169 a_n6641_7124# a_n22897_6995# 0.2797f
C170 a_n7119_7124# a_n22897_6995# 0.2049f
C171 a_n16829_9910# a_n22897_6995# 4.56598f
C172 a_n17107_9910# a_n22897_6995# 2.58447f
C173 a_n22057_9909# a_n22897_6995# 38.1601f
C174 a_n24817_7124# a_n22897_6995# 12.0483f
C175 a_n25295_7124# a_n22897_6995# 0.13378f
C176 a_n14069_7124# a_n22897_6995# 2.82219f
C177 a_n32245_7124# a_n22897_6995# 2.77865f
C178 w_n2704_n7119# a_n22897_6995# 0.2947p
C179 w_n33347_6533# a_n22897_6995# 0.41038p
.ends

