| units: 0.5 tech: gf180mcuD format: MIT
x VREF VSS VCOPY VSUBS s=76800,1520 d=76800,1520 l=282 w=640 x=864 y=-505 nfet_03v3
x a_n2186_n1122# a_n2186_n1122# a_n2186_n1122# VSUBS d=74240,1512 l=282 w=640 x=-1835 y=-505 nfet_03v3
x VREF VSS VCOPY VSUBS s=76800,1520 d=76800,1520 l=282 w=640 x=-475 y=-505 nfet_03v3
x VREF VSS VREF VSUBS s=76800,1520 d=76800,1520 l=282 w=640 x=-1145 y=-505 nfet_03v3
x a_n2186_n1122# a_n2186_n1122# a_n2186_n1122# VSUBS d=74240,1512 l=282 w=640 x=1554 y=-505 nfet_03v3
x VREF VSS VREF VSUBS s=76800,1520 d=76800,1520 l=282 w=640 x=194 y=-505 nfet_03v3
C a_n2186_n1122# VB 0.0
C a_n2186_n1122# VCOPY 1.2
C VCOPY VB 0.0
C VSS VREF 4.6
C a_n2186_n1122# VREF 1.3
C VREF VB 0.0
C VREF VCOPY 0.4
C VSS a_n2186_n1122# 0.5
C VSS VB 0.0
C VSS VCOPY 2.5
C VB0 0.0
C VCOPY0 0.8
R VCOPY 89
C VSS0 1.6
R VSS 192
C VREF0 4.8
R VREF 260
C a_n2186_n1122#0 7.8
R a_n2186_n1122# 1387
