| units: 0.5 tech: gf180mcuD format: MIT
x a_5777_8307# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=5777 y=8687 nfet_03v3
x a_n29950_3049# a_n26898_5979# a_n29950_3049# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-20457 y=5979 pfet_03v3
x a_5777_8307# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6957 y=8687 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5805 y=-7718 nfet_03v3
x a_5657_4411# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6367 y=4411 nfet_03v3
x a_n36440_3049# VSS a_n36440_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-32779 y=543 nfet_03v3
x a_n48062_5772# a_n48182_5979# a_n48062_5772# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-46481 y=5979 pfet_03v3
x a_n48062_5772# a_n48182_5979# a_n48062_5772# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-44111 y=5979 pfet_03v3
x a_n48182_5979# w_n49368_5436# a_n40012_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-39891 y=8885 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=7611 y=-1654 nfet_03v3
x a_5657_4411# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7547 y=4411 nfet_03v3
x a_n1505_n5930# VDD a_n715_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-594 y=-1233 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2192 y=-1233 pfet_03v3
x a_n29950_3049# a_n26898_5979# a_n29950_3049# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-25197 y=5979 pfet_03v3
x a_n36440_3049# VSS a_n30270_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-30149 y=543 nfet_03v3
x a_n39492_5979# a_n36440_3049# a_n39492_5979# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-35139 y=3049 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1793 y=-1233 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5169 y=4411 nfet_03v3
x a_n39492_5979# a_n36440_3049# a_n39492_5979# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-36319 y=3049 nfet_03v3
x VIN a_n715_n5930# a_n195_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-594 y=-5929 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2192 y=-5929 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=7611 y=-7718 nfet_03v3
x a_n36440_3049# VSS a_n36440_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-35139 y=543 nfet_03v3
x a_n29950_3049# a_n26898_5979# a_n29950_3049# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-24407 y=5979 pfet_03v3
x a_n29950_3049# a_n26898_5979# a_n29950_3049# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-26777 y=5979 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1793 y=-5929 pfet_03v3
x a_n1505_n5930# VDD a_75_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=195 y=-1233 pfet_03v3
x a_595_n5930# a_6293_483# a_595_n5930# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6413 y=483 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8155 y=4411 nfet_03v3
x a_n36440_3049# VSS a_n36440_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-31009 y=543 nfet_03v3
x VAUX a_5777_8307# a_1385_n5930# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6367 y=8687 nfet_03v3
x VAUX a_5777_8307# a_1385_n5930# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7547 y=8687 nfet_03v3
x VIN a_75_n5930# a_595_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=195 y=-5929 pfet_03v3
x EN VDD a_n1505_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-199 y=3567 pfet_03v3
x a_n48182_5979# w_n49368_5436# a_n48182_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-42531 y=8885 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5169 y=8687 nfet_03v3
x a_n39492_5979# a_n30270_3049# a_n29950_3049# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-30149 y=3049 nfet_03v3
x a_n26898_5979# w_n49368_5436# a_n26898_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-21247 y=8885 pfet_03v3
x a_6293_483# VSS a_6883_483# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7003 y=-1654 nfet_03v3
x a_n36440_3049# VSS a_n36440_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-33369 y=543 nfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=232000,4232 l=400 w=2000 x=-39083 y=5979 pfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=232000,4232 l=400 w=2000 x=-27585 y=8885 pfet_03v3
x a_1385_n5930# VSS a_5777_8307# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=5777 y=6549 nfet_03v3
x a_n48182_5979# w_n49368_5436# a_n48182_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-47271 y=8885 pfet_03v3
x a_n48062_5772# a_n48182_5979# a_n48062_5772# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-40951 y=5979 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8155 y=8687 nfet_03v3
x a_n26898_5979# w_n49368_5436# a_n26898_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-22827 y=8885 pfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=231884,4230 l=400 w=1999 x=-48869 y=12584 pfet_03v3
x a_1385_n5930# VSS a_5777_8307# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6957 y=6549 nfet_03v3
x a_n29950_3049# a_n18728_5979# a_n18208_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-18607 y=5979 pfet_03v3
x a_n195_n5930# VSS VOUT_VCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7003 y=-7718 nfet_03v3
x a_n48062_5772# a_n48182_5979# a_n48062_5772# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-45691 y=5979 pfet_03v3
x a_n48062_5772# a_n48182_5979# a_n48062_5772# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-43321 y=5979 pfet_03v3
x a_595_n5930# a_6883_483# VOUT_SBCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7003 y=483 nfet_03v3
x VSS VSS VSS VSS d=185600,3432 l=200 w=1600 x=-29541 y=543 nfet_03v3
x a_n36440_3049# VSS a_n36440_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-31599 y=543 nfet_03v3
x a_n48062_12376# a_n26898_12584# a_n26898_5979# w_n49368_5436# s=239880,4238 d=239880,4238 l=400 w=1999 x=-26777 y=12584 pfet_03v3
x VSS VSS VSS VSS d=185600,3432 l=200 w=1600 x=-36927 y=543 nfet_03v3
x a_n29950_3049# a_n26898_5979# a_n29950_3049# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-22037 y=5979 pfet_03v3
x a_n48062_12376# a_n48182_12584# a_n48182_5979# w_n49368_5436# s=239880,4238 d=239880,4238 l=400 w=1999 x=-48061 y=12584 pfet_03v3
x a_n48062_5772# a_n48182_5979# a_n48062_5772# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-44901 y=5979 pfet_03v3
x a_n29950_3049# a_n26898_5979# a_n29950_3049# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-19667 y=5979 pfet_03v3
x a_n48062_5772# a_n48182_5979# a_n48062_5772# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-48061 y=5979 pfet_03v3
x a_n29950_3049# a_n26898_5979# a_n29950_3049# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-23617 y=5979 pfet_03v3
x a_n29950_3049# a_n26898_5979# a_n29950_3049# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-25987 y=5979 pfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=232000,4232 l=400 w=2000 x=-48869 y=5979 pfet_03v3
x a_1385_n5930# VSS a_5657_4411# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6367 y=6549 nfet_03v3
x a_1385_n5930# VSS a_5657_4411# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7547 y=6549 nfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=232000,4232 l=400 w=2000 x=-17799 y=8885 pfet_03v3
x a_n48182_5979# w_n49368_5436# a_n48182_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-41741 y=8885 pfet_03v3
x VSS VSS VSS VSS d=185716,3434 l=200 w=1601 x=-29541 y=3049 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5169 y=6549 nfet_03v3
x a_n48062_5772# a_n40012_5979# a_n39492_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-39891 y=5979 pfet_03v3
x a_n26898_5979# w_n49368_5436# a_n26898_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-20457 y=8885 pfet_03v3
x EN VDD a_n1505_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-989 y=3567 pfet_03v3
x a_n1505_n5930# VDD a_n1505_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1384 y=-1233 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8155 y=6549 nfet_03v3
x a_n36440_3049# VSS a_n36440_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-32189 y=543 nfet_03v3
x a_n48182_5979# w_n49368_5436# a_n48182_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-46481 y=8885 pfet_03v3
x a_n36440_3049# VSS a_n36440_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-35729 y=543 nfet_03v3
x a_n31010_3002# a_n36440_3049# a_n39492_5979# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-31009 y=3049 nfet_03v3
x a_n48182_5979# w_n49368_5436# a_n48182_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-44111 y=8885 pfet_03v3
x VIN a_n1505_n5930# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1384 y=-5929 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1398 y=3567 pfet_03v3
x EN VDD a_n1505_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=590 y=3567 pfet_03v3
x a_n26898_5979# w_n49368_5436# a_n26898_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-25197 y=8885 pfet_03v3
x a_n1505_n5930# VDD a_865_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=985 y=-1233 pfet_03v3
x a_n48062_5772# a_n48182_5979# a_n48062_5772# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-42531 y=5979 pfet_03v3
x a_n26898_5979# w_n49368_5436# a_n26898_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-26777 y=8885 pfet_03v3
x a_6293_483# VSS a_6293_483# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6413 y=-1654 nfet_03v3
x a_n26898_5979# w_n49368_5436# a_n26898_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-24407 y=8885 pfet_03v3
x a_n39492_5979# a_n36440_3049# a_n39492_5979# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-31599 y=3049 nfet_03v3
x a_n29950_3049# a_n26898_5979# a_n29950_3049# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-21247 y=5979 pfet_03v3
x VIN a_865_n5930# a_1385_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=985 y=-5929 pfet_03v3
x a_n39492_5979# a_n36440_3049# a_n39492_5979# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-32779 y=3049 nfet_03v3
x a_n36440_3049# VSS a_n36440_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-33959 y=543 nfet_03v3
x a_n39492_5979# a_n36440_3049# a_n39492_5979# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-33959 y=3049 nfet_03v3
x a_n195_n5930# VSS a_n195_n5930# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6413 y=-7718 nfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=232000,4232 l=400 w=2000 x=-27585 y=5979 pfet_03v3
x a_n48062_5772# a_n48182_5979# a_n48062_5772# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-47271 y=5979 pfet_03v3
x a_n29950_3049# a_n26898_5979# a_n29950_3049# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-22827 y=5979 pfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=232000,4232 l=400 w=2000 x=-39083 y=8885 pfet_03v3
x a_n36440_3049# VSS a_n36440_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-36319 y=543 nfet_03v3
x a_n48182_5979# w_n49368_5436# a_n48182_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-40951 y=8885 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5805 y=483 nfet_03v3
x a_n26898_5979# w_n49368_5436# a_n18728_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-18607 y=8885 pfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=231884,4230 l=400 w=1999 x=-25969 y=12584 pfet_03v3
x VAUX a_5657_4411# VOUT_RCCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=5777 y=4411 nfet_03v3
x a_n39492_5979# a_n36440_3049# a_n39492_5979# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-32189 y=3049 nfet_03v3
x VSS VSS VSS VSS d=185716,3434 l=200 w=1601 x=-36927 y=3049 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-1797 y=3567 pfet_03v3
x VAUX a_5657_4411# VOUT_RCCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6957 y=4411 nfet_03v3
x a_n39492_5979# a_n36440_3049# a_n39492_5979# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-33369 y=3049 nfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=231884,4230 l=400 w=1999 x=-27585 y=12584 pfet_03v3
x a_n48182_5979# w_n49368_5436# a_n48182_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-45691 y=8885 pfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=231884,4230 l=400 w=1999 x=-47253 y=12584 pfet_03v3
x a_n48182_5979# w_n49368_5436# a_n48182_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-43321 y=8885 pfet_03v3
x a_n39492_5979# a_n36440_3049# a_n39492_5979# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-34549 y=3049 nfet_03v3
x a_n36440_3049# VSS a_n36440_3049# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-34549 y=543 nfet_03v3
x a_n39492_5979# a_n36440_3049# a_n39492_5979# VSS s=192120,3442 d=192120,3442 l=200 w=1601 x=-35729 y=3049 nfet_03v3
x a_n26898_5979# w_n49368_5436# a_n26898_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-22037 y=8885 pfet_03v3
x a_n48182_5979# w_n49368_5436# a_n48182_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-44901 y=8885 pfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=232000,4232 l=400 w=2000 x=-17799 y=5979 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=7611 y=483 nfet_03v3
x a_n26898_5979# w_n49368_5436# a_n26898_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-19667 y=8885 pfet_03v3
x a_n48062_5772# a_n48182_5979# a_n48062_5772# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-41741 y=5979 pfet_03v3
x a_n26898_5979# w_n49368_5436# a_n26898_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-25987 y=8885 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5805 y=-1654 nfet_03v3
x a_n48182_5979# w_n49368_5436# a_n48182_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-48061 y=8885 pfet_03v3
x a_n26898_5979# w_n49368_5436# a_n26898_5979# w_n49368_5436# s=240000,4240 d=240000,4240 l=400 w=2000 x=-23617 y=8885 pfet_03v3
x w_n49368_5436# w_n49368_5436# w_n49368_5436# w_n49368_5436# d=232000,4232 l=400 w=2000 x=-48869 y=8885 pfet_03v3
C a_n48062_12376# w_n49368_5436# 5.5
C a_n18208_5979# w_n49368_5436# 1.5
C a_n39492_5979# a_n48062_5772# 0.5
C a_n1505_n5930# VDD 31.5
C a_6883_483# VOUT_SBCM 1.2
C a_n48062_12376# a_n48182_5979# 0.8
C a_n48062_12376# a_n40012_5979# 0.0
C a_5777_8307# a_1385_n5930# 3.0
C a_n715_n5930# a_595_n5930# 0.2
C a_n29950_3049# w_n49368_5436# 15.4
C a_n26898_5979# w_n49368_5436# 47.7
C a_n715_n5930# a_1385_n5930# 0.1
C a_75_n5930# VDD 6.4
C VOUT_RCCM a_1385_n5930# 0.0
C VIN a_n715_n5930# 2.6
C a_n26898_12584# a_n48062_12376# 0.6
C a_n715_n5930# a_n195_n5930# 2.0
C a_n48062_12376# a_n48182_12584# 0.6
C a_n39492_5979# a_n31010_3002# 0.1
C a_595_n5930# VOUT_SBCM 0.2
C VDD a_595_n5930# 1.0
C VDD a_1385_n5930# 2.6
C a_n39492_5979# a_n36440_3049# 36.2
C a_865_n5930# EN 0.2
C a_n26898_12584# a_n26898_5979# 1.0
C VIN VDD 10.3
C a_n48182_5979# w_n49368_5436# 47.7
C a_n40012_5979# w_n49368_5436# 3.1
C a_865_n5930# a_n715_n5930# 0.3
C a_n1505_n5930# a_75_n5930# 1.4
C a_5777_8307# VAUX 3.6
C a_n195_n5930# VDD 1.1
C a_5657_4411# a_1385_n5930# 0.9
C a_6293_483# VOUT_SBCM 0.1
C VOUT_RCCM VAUX 0.6
C a_n48182_5979# a_n40012_5979# 1.0
C a_n26898_12584# w_n49368_5436# 1.4
C a_n48182_12584# w_n49368_5436# 1.4
C a_865_n5930# VDD 5.4
C a_n18208_5979# a_n18728_5979# 0.9
C a_n39492_5979# a_n30270_3049# 0.9
C a_n31010_3002# a_n36440_3049# 0.4
C a_n1505_n5930# a_595_n5930# 0.1
C a_n48182_12584# a_n48182_5979# 1.0
C a_n1505_n5930# a_1385_n5930# 0.8
C a_6883_483# a_595_n5930# 1.5
C a_n39492_5979# a_n29950_3049# 0.3
C VIN a_n1505_n5930# 3.0
C a_n715_n5930# EN 0.0
C a_n18728_5979# a_n29950_3049# 1.0
C VOUT_RCCM a_5777_8307# 0.0
C a_n18728_5979# a_n26898_5979# 1.0
C a_75_n5930# a_595_n5930# 2.0
C a_75_n5930# a_1385_n5930# 0.1
C a_n1505_n5930# a_n195_n5930# 0.1
C VIN a_75_n5930# 0.6
C a_5657_4411# VAUX 3.3
C a_6883_483# a_6293_483# 0.4
C a_75_n5930# a_n195_n5930# 2.0
C a_n39492_5979# w_n49368_5436# 1.8
C a_n48062_5772# w_n49368_5436# 15.1
C a_n31010_3002# a_n30270_3049# 0.0
C a_n18728_5979# w_n49368_5436# 3.1
C VDD EN 7.3
C a_865_n5930# a_n1505_n5930# 2.2
C a_595_n5930# a_1385_n5930# 0.4
C a_n715_n5930# VDD 6.3
C a_n39492_5979# a_n48182_5979# 0.1
C a_n36440_3049# a_n30270_3049# 0.5
C a_n39492_5979# a_n40012_5979# 0.9
C a_n29950_3049# a_n31010_3002# 0.0
C a_n48182_5979# a_n48062_5772# 29.5
C a_n40012_5979# a_n48062_5772# 1.0
C VIN a_595_n5930# 0.6
C VIN a_1385_n5930# 0.6
C a_865_n5930# a_75_n5930# 0.7
C a_n29950_3049# a_n36440_3049# 0.0
C a_n195_n5930# a_595_n5930# 0.5
C a_5777_8307# a_5657_4411# 0.4
C a_n195_n5930# a_1385_n5930# 0.1
C a_6293_483# a_595_n5930# 1.9
C VOUT_RCCM a_5657_4411# 2.2
C VIN a_n195_n5930# 0.6
C a_n195_n5930# VOUT_VCM 0.2
C a_865_n5930# a_595_n5930# 2.0
C a_865_n5930# a_1385_n5930# 2.0
C a_n1505_n5930# EN 1.6
C a_n48062_12376# a_n26898_5979# 0.7
C a_n18208_5979# a_n29950_3049# 0.5
C a_n1505_n5930# a_n715_n5930# 1.7
C a_n18208_5979# a_n26898_5979# 0.1
C a_865_n5930# VIN 0.6
C VAUX a_1385_n5930# 1.7
C a_n29950_3049# a_n30270_3049# 1.1
C a_75_n5930# EN 0.0
C a_865_n5930# a_n195_n5930# 0.1
C a_n715_n5930# a_75_n5930# 0.8
C a_n29950_3049# a_n26898_5979# 29.6
C VOUT_VCM0 3.0
R VOUT_VCM 47
C VOUT_SBCM0 1.7
R VOUT_SBCM 47
C VOUT_RCCM0 3.1
R VOUT_RCCM 107
C VAUX0 16.1
R VAUX 476
C VIN0 2.1
R VIN 414
C EN0 1.4
R EN 198
C VDD0 234.0
R VDD 9009
R VSS 12256
C a_6883_483#0 2.9
R a_6883_483# 107
C a_6293_483#0 6.4
R a_6293_483# 219
C a_5657_4411#0 8.5
R a_5657_4411# 340
C a_5777_8307#0 7.7
R a_5777_8307# 335
C a_1385_n5930#0 12.2
R a_1385_n5930# 486
C a_595_n5930#0 4.5
R a_595_n5930# 291
C a_n195_n5930#0 7.8
R a_n195_n5930# 290
C a_865_n5930#0 0.2
R a_865_n5930# 269
C a_75_n5930#0 0.0
R a_75_n5930# 269
C a_n715_n5930#0 0.0
R a_n715_n5930# 269
C a_n1505_n5930#0 2.7
R a_n1505_n5930# 974
C a_n30270_3049#0 2.8
R a_n30270_3049# 191
C a_n36440_3049#0 40.2
R a_n36440_3049# 2963
C a_n31010_3002#0 0.3
R a_n31010_3002# 62
C a_n18208_5979#0 0.4
R a_n18208_5979# 123
C a_n29950_3049#0 5.4
R a_n29950_3049# 2091
C a_n18728_5979#0 0.3
R a_n18728_5979# 260
C a_n39492_5979#0 13.0
R a_n39492_5979# 1995
C a_n48062_5772#0 2.8
R a_n48062_5772# 1998
C a_n40012_5979#0 0.3
R a_n40012_5979# 260
C a_n26898_5979#0 3.2
R a_n26898_5979# 3505
C a_n26898_12584#0 0.2
R a_n26898_12584# 122
C a_n48182_5979#0 3.2
R a_n48182_5979# 3505
C a_n48182_12584#0 0.2
R a_n48182_12584# 122
C a_n48062_12376#0 6.3
R a_n48062_12376# 122
C w_n49368_5436#0 495.4
R w_n49368_5436# 26599
