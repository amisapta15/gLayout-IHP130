| units: 500000 tech: sky130A format: MIT
x a_n32245_7124# w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-26208 y=9909 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=5351 y=8553 sky130_fd_pr__nfet_01v8
x a_n22057_9909# a_n22897_6995# a_n17107_9910# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-17028 y=7524 sky130_fd_pr__nfet_01v8
x a_200_n5640# a_6260_503# a_200_n5640# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6338 y=503 sky130_fd_pr__nfet_01v8
x VAUX a_n32245_7124# VAUX w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-27532 y=7124 sky130_fd_pr__pfet_01v8
x a_5835_4440# a_5757_4829# VOUT_RCCM a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6759 y=4829 sky130_fd_pr__nfet_01v8
x w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# d=156000,4156 l=400 w=2000 x=1477 y=3681 sky130_fd_pr__pfet_01v8
x EN w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-32166 y=13534 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=7284 y=503 sky130_fd_pr__nfet_01v8
x a_6260_503# a_n22897_6995# a_6722_503# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6800 y=-1359 sky130_fd_pr__nfet_01v8
x a_n22057_9909# a_n22897_6995# a_n22057_9909# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-17820 y=7524 sky130_fd_pr__nfet_01v8
x a_n24817_7124# a_n22057_9909# a_n24817_7124# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-17820 y=9909 sky130_fd_pr__nfet_01v8
x a_n16829_9910# a_n14069_7124# a_n16829_9910# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-8032 y=7124 sky130_fd_pr__pfet_01v8
x a_n16829_9910# a_n14069_7124# a_n16829_9910# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-12004 y=7124 sky130_fd_pr__pfet_01v8
x a_n22057_9909# a_n22897_6995# a_n22057_9909# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-20130 y=7524 sky130_fd_pr__nfet_01v8
x a_n22057_9909# a_n22897_6995# a_n22057_9909# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-21516 y=7524 sky130_fd_pr__nfet_01v8
x a_n24817_7124# a_n22057_9909# a_n24817_7124# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-21516 y=9909 sky130_fd_pr__nfet_01v8
x a_n24817_7124# a_n22057_9909# a_n24817_7124# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-20130 y=9909 sky130_fd_pr__nfet_01v8
x a_5757_4829# a_n22897_6995# a_5835_4440# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=7221 y=4829 sky130_fd_pr__nfet_01v8
x a_n14069_7124# w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-8694 y=9909 sky130_fd_pr__pfet_01v8
x a_n14069_7124# w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-12666 y=9909 sky130_fd_pr__pfet_01v8
x w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# d=156078,4158 l=400 w=2001 x=-2207 y=-5639 sky130_fd_pr__pfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-14674 y=9909 sky130_fd_pr__pfet_01v8
x w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# d=156078,4158 l=400 w=2001 x=1808 y=-5639 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=5351 y=4829 sky130_fd_pr__nfet_01v8
x EN w_n2704_n7119# a_n1602_n5640# w_n2704_n7119# s=156000,4156 d=156000,4156 l=400 w=2000 x=-530 y=3681 sky130_fd_pr__pfet_01v8
x a_n22057_9909# a_n22897_6995# a_n22057_9909# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-18282 y=7524 sky130_fd_pr__nfet_01v8
x a_n22057_9909# a_n22897_6995# a_n22057_9909# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-19668 y=7524 sky130_fd_pr__nfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=7705 y=6691 sky130_fd_pr__nfet_01v8
x a_n16829_9910# a_n14069_7124# a_n16829_9910# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-13990 y=7124 sky130_fd_pr__pfet_01v8
x a_n24817_7124# a_n22057_9909# a_n24817_7124# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-18282 y=9909 sky130_fd_pr__nfet_01v8
x a_n24817_7124# a_n22057_9909# a_n24817_7124# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-19668 y=9909 sky130_fd_pr__nfet_01v8
x a_862_n5640# a_n22897_6995# a_5835_8163# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=5835 y=6691 sky130_fd_pr__nfet_01v8
x EN w_n2704_n7119# a_n1602_n5640# w_n2704_n7119# s=156000,4156 d=156000,4156 l=400 w=2000 x=793 y=3681 sky130_fd_pr__pfet_01v8
x VAUX a_n32245_7124# VAUX w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-26208 y=7124 sky130_fd_pr__pfet_01v8
x a_n462_n5640# a_n22897_6995# VOUT_VCM a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6800 y=-7548 sky130_fd_pr__nfet_01v8
x w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# d=156000,4156 l=400 w=2000 x=1808 y=-992 sky130_fd_pr__pfet_01v8
x a_n14069_7124# w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-10680 y=9909 sky130_fd_pr__pfet_01v8
x a_862_n5640# a_n22897_6995# a_5757_4829# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6297 y=6691 sky130_fd_pr__nfet_01v8
x a_n32245_7124# w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-32166 y=9909 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=124800,3356 l=200 w=1600 x=-16544 y=7524 sky130_fd_pr__nfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-24532 y=7124 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=7705 y=8553 sky130_fd_pr__nfet_01v8
x w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# d=156000,4156 l=400 w=2000 x=-1876 y=3681 sky130_fd_pr__pfet_01v8
x a_5835_8163# a_n22897_6995# a_5835_4440# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=5835 y=8553 sky130_fd_pr__nfet_01v8
x a_n16829_9910# a_n14069_7124# a_n16829_9910# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-8694 y=7124 sky130_fd_pr__pfet_01v8
x a_n16829_9910# a_n14069_7124# a_n16829_9910# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-12666 y=7124 sky130_fd_pr__pfet_01v8
x a_n1602_n5640# w_n2704_n7119# a_n278_n5640# w_n2704_n7119# s=156000,4156 d=156000,4156 l=400 w=2000 x=-199 y=-992 sky130_fd_pr__pfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-6356 y=9910 sky130_fd_pr__pfet_01v8
x a_n32245_7124# w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-28856 y=9909 sky130_fd_pr__pfet_01v8
x a_n1602_n5640# w_n2704_n7119# a_1046_n5640# w_n2704_n7119# s=156000,4156 d=156000,4156 l=400 w=2000 x=1124 y=-992 sky130_fd_pr__pfet_01v8
x a_n32245_7124# w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-28194 y=9909 sky130_fd_pr__pfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-14674 y=7124 sky130_fd_pr__pfet_01v8
x a_n32245_7124# w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-30842 y=9909 sky130_fd_pr__pfet_01v8
x a_n1524_n6691# a_n278_n5640# a_200_n5640# w_n2704_n7119# s=156078,4158 d=156078,4158 l=400 w=2001 x=-199 y=-5639 sky130_fd_pr__pfet_01v8
x a_n32245_7124# w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-30180 y=9909 sky130_fd_pr__pfet_01v8
x a_n1602_n5640# w_n2704_n7119# a_384_n5640# w_n2704_n7119# s=156000,4156 d=156000,4156 l=400 w=2000 x=462 y=-992 sky130_fd_pr__pfet_01v8
x a_5835_4440# a_5835_8163# a_862_n5640# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6297 y=8553 sky130_fd_pr__nfet_01v8
x a_6260_503# a_n22897_6995# a_6260_503# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6338 y=-1359 sky130_fd_pr__nfet_01v8
x a_n16829_9910# a_n7119_7124# a_n6641_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-7040 y=7124 sky130_fd_pr__pfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-32850 y=9909 sky130_fd_pr__pfet_01v8
x a_n14069_7124# w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-9356 y=9909 sky130_fd_pr__pfet_01v8
x a_n14069_7124# w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-13328 y=9909 sky130_fd_pr__pfet_01v8
x a_n22057_9909# a_n22897_6995# a_n22057_9909# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-19206 y=7524 sky130_fd_pr__nfet_01v8
x a_n24817_7124# a_n22057_9909# a_n24817_7124# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-19206 y=9909 sky130_fd_pr__nfet_01v8
x EN w_n2704_n7119# a_n1602_n5640# w_n2704_n7119# s=156000,4156 d=156000,4156 l=400 w=2000 x=-1192 y=3681 sky130_fd_pr__pfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-32850 y=13534 sky130_fd_pr__pfet_01v8
x a_n16829_9910# a_n14069_7124# a_n16829_9910# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-10680 y=7124 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=7284 y=-1359 sky130_fd_pr__nfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=7705 y=4829 sky130_fd_pr__nfet_01v8
x a_n32245_7124# w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-26870 y=9909 sky130_fd_pr__pfet_01v8
x a_n1524_n6691# a_1046_n5640# VOUT_VIN w_n2704_n7119# s=156078,4158 d=156078,4158 l=400 w=2001 x=1124 y=-5639 sky130_fd_pr__pfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-14674 y=13534 sky130_fd_pr__pfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-31482 y=13534 sky130_fd_pr__pfet_01v8
x VAUX a_n32245_7124# VAUX w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-32166 y=7124 sky130_fd_pr__pfet_01v8
x VAUX a_n25295_7124# a_n24817_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-25216 y=7124 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=5854 y=503 sky130_fd_pr__nfet_01v8
x a_5835_4440# a_5757_4829# VOUT_RCCM a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=5835 y=4829 sky130_fd_pr__nfet_01v8
x a_n462_n5640# a_n22897_6995# a_n462_n5640# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6338 y=-7548 sky130_fd_pr__nfet_01v8
x a_n14069_7124# w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-11342 y=9909 sky130_fd_pr__pfet_01v8
x a_5757_4829# a_n22897_6995# a_5835_4440# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6297 y=4829 sky130_fd_pr__nfet_01v8
x VAUX a_n32245_7124# VAUX w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-28856 y=7124 sky130_fd_pr__pfet_01v8
x a_n1524_n6691# a_n1602_n5640# a_n1524_n6691# w_n2704_n7119# s=156078,4158 d=156078,4158 l=400 w=2001 x=-1523 y=-5639 sky130_fd_pr__pfet_01v8
x a_n1602_n5640# w_n2704_n7119# a_n940_n5640# w_n2704_n7119# s=156000,4156 d=156000,4156 l=400 w=2000 x=-861 y=-992 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=7284 y=-7548 sky130_fd_pr__nfet_01v8
x VAUX a_n32245_7124# VAUX w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-28194 y=7124 sky130_fd_pr__pfet_01v8
x VAUX a_n32245_7124# VAUX w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-30842 y=7124 sky130_fd_pr__pfet_01v8
x a_n22057_9909# a_n22897_6995# a_n22057_9909# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-18744 y=7524 sky130_fd_pr__nfet_01v8
x VAUX a_n32245_7124# VAUX w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-30180 y=7124 sky130_fd_pr__pfet_01v8
x a_n1602_n5640# w_n2704_n7119# a_n1602_n5640# w_n2704_n7119# s=156000,4156 d=156000,4156 l=400 w=2000 x=-1523 y=-992 sky130_fd_pr__pfet_01v8
x a_n24817_7124# a_n22057_9909# a_n24817_7124# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-18744 y=9909 sky130_fd_pr__nfet_01v8
x a_n22057_9909# a_n22897_6995# a_n22057_9909# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-21054 y=7524 sky130_fd_pr__nfet_01v8
x a_n24817_7124# a_n17107_9910# a_n16829_9910# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-17028 y=9910 sky130_fd_pr__nfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-32850 y=7124 sky130_fd_pr__pfet_01v8
x a_n24817_7124# a_n22057_9909# a_n24817_7124# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-21054 y=9909 sky130_fd_pr__nfet_01v8
x a_n16829_9910# a_n14069_7124# a_n16829_9910# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-9356 y=7124 sky130_fd_pr__pfet_01v8
x a_n16829_9910# a_n14069_7124# a_n16829_9910# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-13328 y=7124 sky130_fd_pr__pfet_01v8
x a_n32245_7124# w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-29518 y=9909 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=5854 y=-1359 sky130_fd_pr__nfet_01v8
x a_n32245_7124# w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-31504 y=9909 sky130_fd_pr__pfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-24532 y=9910 sky130_fd_pr__pfet_01v8
x VAUX a_n32245_7124# VAUX w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-26870 y=7124 sky130_fd_pr__pfet_01v8
x a_862_n5640# a_n22897_6995# a_5835_8163# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6759 y=6691 sky130_fd_pr__nfet_01v8
x a_n14069_7124# w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-10018 y=9909 sky130_fd_pr__pfet_01v8
x a_n16829_9910# a_n14069_7124# a_n16829_9910# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-11342 y=7124 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=124800,3356 l=200 w=1600 x=-22462 y=7524 sky130_fd_pr__nfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=124800,3356 l=200 w=1600 x=-22462 y=9909 sky130_fd_pr__nfet_01v8
x a_862_n5640# a_n22897_6995# a_5757_4829# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=7221 y=6691 sky130_fd_pr__nfet_01v8
x a_n32245_7124# w_n33347_6533# a_n32245_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-27532 y=9909 sky130_fd_pr__pfet_01v8
x a_n14069_7124# w_n33347_6533# a_n7119_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-7040 y=9910 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=5854 y=-7548 sky130_fd_pr__nfet_01v8
x a_n22057_9909# a_n22897_6995# a_n22057_9909# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-20592 y=7524 sky130_fd_pr__nfet_01v8
x a_n22057_9909# a_n22897_6995# a_n22057_9909# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-21978 y=7524 sky130_fd_pr__nfet_01v8
x a_n24817_7124# a_n22057_9909# a_n24817_7124# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-21978 y=9909 sky130_fd_pr__nfet_01v8
x a_n24817_7124# a_n22057_9909# a_n24817_7124# a_n22897_6995# s=124800,3356 d=124800,3356 l=200 w=1600 x=-20592 y=9909 sky130_fd_pr__nfet_01v8
x a_200_n5640# a_6722_503# VOUT_SBCM a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6800 y=503 sky130_fd_pr__nfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=62400,1756 l=200 w=800 x=5351 y=6691 sky130_fd_pr__nfet_01v8
x w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# d=156000,4156 l=400 w=2000 x=-2207 y=-992 sky130_fd_pr__pfet_01v8
x a_5835_8163# a_n22897_6995# a_5835_4440# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=6759 y=8553 sky130_fd_pr__nfet_01v8
x a_n1524_n6691# a_n940_n5640# a_n462_n5640# w_n2704_n7119# s=156078,4158 d=156078,4158 l=400 w=2001 x=-861 y=-5639 sky130_fd_pr__pfet_01v8
x a_n14069_7124# w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-8032 y=9909 sky130_fd_pr__pfet_01v8
x a_n14069_7124# w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-12004 y=9909 sky130_fd_pr__pfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-13306 y=13534 sky130_fd_pr__pfet_01v8
x VAUX a_n32245_7124# VAUX w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-29518 y=7124 sky130_fd_pr__pfet_01v8
x a_n32245_7124# w_n33347_6533# a_n25295_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-25216 y=9910 sky130_fd_pr__pfet_01v8
x a_n14069_7124# w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-13990 y=9909 sky130_fd_pr__pfet_01v8
x a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# d=124800,3356 l=200 w=1600 x=-16544 y=9910 sky130_fd_pr__nfet_01v8
x VAUX a_n32245_7124# VAUX w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-31504 y=7124 sky130_fd_pr__pfet_01v8
x a_5835_4440# a_5835_8163# a_862_n5640# a_n22897_6995# s=62400,1756 d=62400,1756 l=200 w=800 x=7221 y=8553 sky130_fd_pr__nfet_01v8
x w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# d=156000,4156 l=400 w=2000 x=-6356 y=7124 sky130_fd_pr__pfet_01v8
x a_n1524_n6691# a_384_n5640# a_862_n5640# w_n2704_n7119# s=156078,4158 d=156078,4158 l=400 w=2001 x=462 y=-5639 sky130_fd_pr__pfet_01v8
x EN w_n33347_6533# a_n14069_7124# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-13990 y=13534 sky130_fd_pr__pfet_01v8
x EN w_n2704_n7119# a_n1602_n5640# w_n2704_n7119# s=156000,4156 d=156000,4156 l=400 w=2000 x=131 y=3681 sky130_fd_pr__pfet_01v8
x a_n16829_9910# a_n14069_7124# a_n16829_9910# w_n33347_6533# s=156000,4156 d=156000,4156 l=400 w=2000 x=-10018 y=7124 sky130_fd_pr__pfet_01v8
C VAUX li_9462_n10101# 0.0
C a_n16829_9910# a_n24817_7124# 0.5
C VOUT_RCCM li_9462_n10101# 0.1
C VOUT_VIN a_5835_4440# 0.1
C w_n2704_n7119# a_1046_n5640# 5.8
C a_5757_4829# VOUT_RCCM 1.8
C a_1046_n5640# a_384_n5640# 0.6
C a_n940_n5640# EN 0.0
C a_n16829_9910# a_n17107_9910# 0.9
C a_6260_503# a_6722_503# 0.4
C a_n1524_n6691# a_200_n5640# 0.9
C a_n25295_7124# a_n32245_7124# 1.4
C a_n940_n5640# a_862_n5640# 0.1
C a_n278_n5640# a_200_n5640# 2.4
C li_n5290_9325# a_5835_4440# 0.0
C a_862_n5640# a_n462_n5640# 0.1
C a_n7119_7124# a_n14069_7124# 1.4
C a_n25295_7124# a_n24817_7124# 0.8
C a_n16829_9910# w_n2704_n7119# 0.0
C a_n16829_9910# w_n33347_6533# 14.7
C EN a_n25295_7124# 0.0
C a_n940_n5640# w_n2704_n7119# 6.6
C a_200_n5640# a_1046_n5640# 0.1
C VOUT_VIN li_n5290_9325# 0.1
C a_n940_n5640# a_384_n5640# 0.3
C a_n6641_7124# li_n5290_9325# 0.0
C w_n2704_n7119# a_n462_n5640# 1.1
C EN a_n7119_7124# 0.0
C VOUT_VIN a_n1524_n6691# 0.8
C a_200_n5640# VOUT_SBCM 0.3
C VOUT_VIN a_n278_n5640# 0.1
C a_n462_n5640# a_384_n5640# 0.1
C li_n32467_15897# VDD 0.1
C a_n25295_7124# VAUX 1.2
C a_5757_4829# a_5835_4440# 3.3
C a_n25295_7124# w_n33347_6533# 2.9
C VOUT_VIN li_9462_n10101# 0.1
C VOUT_VIN a_1046_n5640# 2.4
C EN a_n1602_n5640# 3.2
C a_n940_n5640# a_200_n5640# 0.1
C li_n32467_15897# a_n32245_7124# 0.0
C a_n7119_7124# w_n33347_6533# 2.9
C a_n1602_n5640# a_862_n5640# 0.4
C a_n1524_n6691# a_n278_n5640# 0.9
C a_200_n5640# a_n462_n5640# 0.7
C a_n24817_7124# a_n32245_7124# 0.1
C EN a_n32245_7124# 1.2
C EN a_n14069_7124# 1.2
C a_n1524_n6691# li_n3142_n10147# 0.0
C li_n32467_15897# EN 0.0
C a_n1602_n5640# w_n2704_n7119# 43.9
C li_6128_10166# a_5835_8163# 0.0
C a_n6641_7124# a_n16829_9910# 0.8
C a_n1524_n6691# a_1046_n5640# 0.9
C a_n278_n5640# a_1046_n5640# 0.3
C a_862_n5640# a_5835_8163# 2.8
C a_n1602_n5640# a_384_n5640# 2.0
C VOUT_VIN a_n940_n5640# 0.1
C VAUX a_n32245_7124# 30.7
C EN li_6128_10166# 0.8
C a_n17107_9910# a_n24817_7124# 1.0
C a_6722_503# a_200_n5640# 1.3
C li_n32467_15897# VAUX 0.5
C VOUT_VIN a_n462_n5640# 0.1
C a_n32245_7124# w_n33347_6533# 48.7
C a_n14069_7124# w_n33347_6533# 48.7
C li_n32467_15897# w_n33347_6533# 1.1
C VAUX a_n24817_7124# 0.8
C a_5835_8163# VOUT_RCCM 0.0
C EN VAUX 0.0
C a_n24817_7124# w_n33347_6533# 1.7
C li_6128_10166# VAUX 0.5
C li_9462_n10101# VOUT_SBCM 0.1
C a_6260_503# a_200_n5640# 1.8
C EN w_n2704_n7119# 13.8
C a_n1602_n5640# a_200_n5640# 0.1
C EN w_n33347_6533# 6.8
C a_n940_n5640# a_n1524_n6691# 2.7
C a_n940_n5640# a_n278_n5640# 0.7
C a_862_n5640# VOUT_RCCM 0.0
C a_862_n5640# w_n2704_n7119# 1.7
C EN a_384_n5640# 0.0
C li_n3142_n10147# li_9474_n10147# 0.0
C a_n6641_7124# a_n7119_7124# 0.8
C a_n17107_9910# w_n33347_6533# 0.0
C VIN li_9462_n10101# 0.0
C a_n1524_n6691# a_n462_n5640# 0.9
C a_862_n5640# a_384_n5640# 2.3
C li_9474_n10147# li_9462_n10101# 0.0
C a_n278_n5640# a_n462_n5640# 1.9
C a_n22057_9909# a_n24817_7124# 36.2
C w_n2704_n7119# VAUX 0.0
C VAUX w_n33347_6533# 15.1
C a_n940_n5640# a_1046_n5640# 0.3
C w_n2704_n7119# w_n33347_6533# 4.7
C li_n5290_9325# a_n7119_7124# 0.0
C li_6128_10166# VSS 0.1
C w_n2704_n7119# a_384_n5640# 6.7
C VOUT_VIN a_n1602_n5640# 0.6
C a_n17107_9910# a_n22057_9909# 0.7
C a_n462_n5640# a_1046_n5640# 0.1
C a_200_n5640# a_862_n5640# 0.3
C a_5835_8163# a_5835_4440# 3.6
C VOUT_VCM li_9462_n10101# 0.1
C a_n6641_7124# a_n14069_7124# 0.0
C li_6128_10166# a_5835_4440# 0.0
C a_862_n5640# a_5835_4440# 1.5
C VOUT_VIN a_5835_8163# 0.0
C a_200_n5640# w_n2704_n7119# 1.0
C a_n1524_n6691# a_n1602_n5640# 3.8
C a_n278_n5640# a_n1602_n5640# 2.0
C a_200_n5640# a_384_n5640# 1.9
C a_n940_n5640# a_n462_n5640# 2.4
C VOUT_VIN li_6128_10166# 0.8
C VOUT_VIN a_862_n5640# 3.0
C a_6722_503# VOUT_SBCM 1.0
C a_5835_4440# VOUT_RCCM 0.7
C a_n1602_n5640# a_1046_n5640# 2.7
C a_n7119_7124# a_n16829_9910# 1.2
C EN li_n5290_9325# 0.0
C a_6260_503# VOUT_SBCM 0.1
C VOUT_VIN w_n2704_n7119# 2.6
C li_n5290_9325# a_862_n5640# 0.1
C VOUT_VCM a_n462_n5640# 0.3
C a_n6641_7124# w_n33347_6533# 1.4
C EN a_n278_n5640# 0.0
C VOUT_VIN a_384_n5640# 0.1
C a_n1524_n6691# a_862_n5640# 0.9
C a_n278_n5640# a_862_n5640# 0.1
C a_5835_8163# a_5757_4829# 0.3
C EN li_9462_n10101# 0.1
C li_n5290_9325# w_n33347_6533# 0.0
C a_n940_n5640# a_n1602_n5640# 2.3
C EN a_1046_n5640# 0.2
C a_n1524_n6691# w_n2704_n7119# 14.3
C a_n278_n5640# w_n2704_n7119# 6.6
C a_862_n5640# a_1046_n5640# 1.9
C a_862_n5640# a_5757_4829# 1.1
C a_n16829_9910# a_n14069_7124# 30.7
C a_n1602_n5640# a_n462_n5640# 0.1
C a_n1524_n6691# a_384_n5640# 0.9
C VOUT_VIN a_200_n5640# 0.1
C a_n278_n5640# a_384_n5640# 0.7
C VIN0 0.1
R VIN 13
C VSS0 0.1
R VSS 25
C VDD0 0.1
R VDD 23
C VOUT_VCM0 5.5
R VOUT_VCM 1547
C VOUT_VIN0 10.2
R VOUT_VIN 5813
C VOUT_SBCM0 4.2
R VOUT_SBCM 1547
C VOUT_RCCM0 5.3
R VOUT_RCCM 3305
C VAUX0 25.3
R VAUX 64244
C EN0 22.9
R EN 4333
C li_9474_n10147#0 0.0
R li_9474_n10147# 13
C li_n3142_n10147#0 5.8
R li_n3142_n10147# 2786
C li_n5290_9325#0 4.6
R li_n5290_9325# 2221
C li_9462_n10101#0 18.9
R li_9462_n10101# 9079
C li_6128_10166#0 41.1
R li_6128_10166# 383
C li_n32467_15897#0 92.1
R li_n32467_15897# 884
C a_n462_n5640#0 7.9
R a_n462_n5640# 8073
C a_n1524_n6691#0 4.1
R a_n1524_n6691# 10567
C a_6722_503#0 2.6
R a_6722_503# 3248
C a_6260_503#0 6.1
R a_6260_503# 4045
C a_200_n5640#0 5.0
R a_200_n5640# 8075
C a_1046_n5640#0 0.0
R a_1046_n5640# 11851
R a_384_n5640# 11847
R a_n278_n5640# 11847
R a_n940_n5640# 11847
C a_5757_4829#0 7.6
R a_5757_4829# 7573
C a_n1602_n5640#0 2.2
R a_n1602_n5640# 39933
C a_862_n5640#0 12.0
R a_862_n5640# 10760
C a_5835_4440#0 11.7
R a_5835_4440# 8525
C a_5835_8163#0 6.9
R a_5835_8163# 7549
C a_n6641_7124#0 0.3
R a_n6641_7124# 5508
C a_n7119_7124#0 0.2
R a_n7119_7124# 11384
C a_n16829_9910#0 4.6
R a_n16829_9910# 66999
C a_n17107_9910#0 2.6
R a_n17107_9910# 5889
C a_n22057_9909#0 38.2
R a_n22057_9909# 67839
C a_n24817_7124#0 12.0
R a_n24817_7124# 42550
C a_n25295_7124#0 0.1
R a_n25295_7124# 11384
C a_n14069_7124#0 2.8
R a_n14069_7124# 129057
C a_n32245_7124#0 2.8
R a_n32245_7124# 129057
C w_n2704_n7119#0 294.7
R w_n2704_n7119# 178123
C w_n33347_6533#0 410.4
R w_n33347_6533# 411406
R a_n22897_6995# 280823
