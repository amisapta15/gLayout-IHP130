* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu9t5v0__tieh$2 VDD VSS Z VNW VPW a_125_157#
X0 Z a_125_157# VDD VNW pfet_05v0 ad=0.396p pd=2.68u as=0.396p ps=2.68u w=0.9u l=0.5u
X1 a_125_157# a_125_157# VSS VPW nfet_05v0 ad=0.2904p pd=2.2u as=0.2904p ps=2.2u w=0.66u l=0.6u
C0 VDD Z 0.05696f
C1 VSS a_125_157# 0.05594f
C2 VDD VSS 0.02071f
C3 VNW a_125_157# 0.13984f
C4 VNW VDD 0.13685f
C5 VDD a_125_157# 0.02505f
C6 VNW Z 0.01694f
C7 Z a_125_157# 0.0165f
C8 VNW VSS 0.01055f
C9 VSS VPW 0.31582f
C10 Z VPW 0.02933f
C11 VDD VPW 0.23581f
C12 VNW VPW 1.19226f
C13 a_125_157# VPW 0.37323f
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__tiel$3 VDD VSS ZN VNW VPW a_124_157#
X0 ZN a_124_157# VSS VPW nfet_05v0 ad=0.2904p pd=2.2u as=0.2904p ps=2.2u w=0.66u l=0.6u
X1 a_124_157# a_124_157# VDD VNW pfet_05v0 ad=0.396p pd=2.68u as=0.396p ps=2.68u w=0.9u l=0.5u
C0 VDD VSS 0.02032f
C1 ZN a_124_157# 0.02544f
C2 VDD ZN 0
C3 VNW a_124_157# 0.15591f
C4 VSS ZN 0.03448f
C5 VNW VDD 0.13657f
C6 VDD a_124_157# 0.08266f
C7 VNW VSS 0.01117f
C8 VSS a_124_157# 0.03129f
C9 VNW ZN 0
C10 ZN VPW 0.02686f
C11 VSS VPW 0.31286f
C12 VDD VPW 0.23555f
C13 VNW VPW 1.19226f
C14 a_124_157# VPW 0.3723f
.ends

.subckt sc_tieh_tiel$1 tieH tieL gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# VDD
+ gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# VSS
Xgf180mcu_fd_sc_mcu9t5v0__tieh$2_0 VDD VSS tieH VDD VSS gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157#
+ gf180mcu_fd_sc_mcu9t5v0__tieh$2
Xgf180mcu_fd_sc_mcu9t5v0__tiel$3_0 VDD VSS tieL VDD VSS gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157#
+ gf180mcu_fd_sc_mcu9t5v0__tiel$3
C0 tieH VSS 0.01457f
C1 gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# VDD 0.02329f
C2 gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# VDD 0.00888f
C3 gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# tieL 0.01483f
C4 VDD VSS 0.29762f
C5 gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# tieL 0
C6 tieL VSS 0.08309f
C7 gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# 0.0027f
C8 tieH VDD 0.08219f
C9 gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# VSS 0.01505f
C10 tieH tieL 0.01031f
C11 gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# VSS 0.02873f
C12 tieL VDD 0.03191f
C13 tieH gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# 0.00414f
C14 VSS 0 1.29627f
C15 VDD 0 3.38527f
C16 tieL 0 0.16778f
C17 gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# 0 0.3723f
C18 tieH 0 0.13137f
C19 gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# 0 0.37323f
.ends

.subckt ppolyf_u_9H3LNU$2 a_n224793_504053# w_n225009_503837# a_n224793_506155# VSUBS
X0 a_n224793_506155# a_n224793_504053# w_n225009_503837# ppolyf_u r_width=40u r_length=10u
C0 a_n224793_504053# w_n225009_503837# 6.29946f
C1 a_n224793_506155# w_n225009_503837# 6.29946f
C2 a_n224793_504053# VSUBS 4.5322f
C3 a_n224793_506155# VSUBS 4.5322f
C4 w_n225009_503837# VSUBS 72.7085f
.ends

.subckt diode_nd2ps_06v0_MV3SZ3$2 a_505271_219793# a_503039_219793# a_507503_219793#
+ a_500807_219793# a_500655_219641#
D0 a_500655_219641# a_505271_219793# diode_nd2ps_06v0 pj=40u area=99.99999p
D1 a_500655_219641# a_500807_219793# diode_nd2ps_06v0 pj=40u area=99.99999p
D2 a_500655_219641# a_503039_219793# diode_nd2ps_06v0 pj=40u area=99.99999p
D3 a_500655_219641# a_507503_219793# diode_nd2ps_06v0 pj=40u area=99.99999p
C0 a_507503_219793# a_500655_219641# 3.83321f
C1 a_505271_219793# a_500655_219641# 3.83321f
C2 a_503039_219793# a_500655_219641# 3.83321f
C3 a_500807_219793# a_500655_219641# 3.83321f
.ends

.subckt diode_pd2nw_06v0_5DG9HC$2 a_507479_219793# a_500831_219793# w_500655_219617#
+ a_503047_219793# a_505263_219793# a_500511_219473#
D0 a_500831_219793# w_500655_219617# diode_pd2nw_06v0 pj=40u area=99.99999p
D1 a_507479_219793# w_500655_219617# diode_pd2nw_06v0 pj=40u area=99.99999p
D2 a_503047_219793# w_500655_219617# diode_pd2nw_06v0 pj=40u area=99.99999p
D3 a_505263_219793# w_500655_219617# diode_pd2nw_06v0 pj=40u area=99.99999p
C0 w_500655_219617# a_503047_219793# 4.17112f
C1 a_505263_219793# w_500655_219617# 4.17112f
C2 a_500831_219793# w_500655_219617# 4.17112f
C3 a_507479_219793# w_500655_219617# 4.17112f
C4 w_500655_219617# a_500511_219473# 73.4915f
.ends

.subckt io_secondary_5p0$1 m1_512035_219553# m1_499212_228525# VSUBS m1_497955_232243#
Xppolyf_u_9H3LNU_0 m1_499212_228525# m1_497955_232243# m1_512035_219553# VSUBS ppolyf_u_9H3LNU$2
Xdiode_nd2ps_06v0_MV3SZ3_0 m1_499212_228525# m1_499212_228525# m1_499212_228525# m1_499212_228525#
+ VSUBS diode_nd2ps_06v0_MV3SZ3$2
Xdiode_pd2nw_06v0_5DG9HC_0 m1_499212_228525# m1_499212_228525# m1_497955_232243# m1_499212_228525#
+ m1_499212_228525# VSUBS diode_pd2nw_06v0_5DG9HC$2
C0 m1_499212_228525# m1_497955_232243# 16.86721f
C1 m1_512035_219553# m1_497955_232243# 11.99056f
C2 m1_499212_228525# VSUBS 0.15225p
C3 m1_512035_219553# VSUBS 5.38418f
C4 m1_497955_232243# VSUBS 0.17048p
.ends

.subckt M a_402461_244568# a_410134_251737# a_408568_255933# a_403521_244568# a_365828_259091#
+ a_411044_251737# a_409618_256263# a_409618_260539# a_404831_244568# a_401271_243528#
+ a_409818_256643# a_403251_244568# a_365828_265695# a_404311_244568# a_376520_259212#
+ a_401941_244568# a_395682_259299# a_404041_244568# a_409498_256643# a_402731_244568#
+ a_401151_244568# a_411044_242557# w_364522_258756#
X0 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0.4068n ps=1.46136m w=10u l=2u
X1 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X2 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X3 a_402461_244568# a_401271_243528# a_401941_244568# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X4 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X5 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X6 a_404311_244568# a_401151_244568# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X7 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X8 a_374398_259299# a_365828_259091# a_373878_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X9 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X10 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X11 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X12 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X13 a_401151_244568# a_401151_244568# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X14 a_404041_244568# a_409618_256263# a_409618_260539# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X15 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.64p pd=17.16u as=0.1744n ps=0.65672m w=8u l=1u
X16 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X17 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X18 a_409618_256263# a_409618_260539# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X19 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X20 a_409618_256263# a_409498_256643# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X21 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X22 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X23 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X24 a_409618_256263# a_409618_260539# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X25 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X26 a_401151_244568# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X27 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X28 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X29 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X30 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X31 a_401151_244568# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X32 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X33 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X34 a_404041_244568# a_401271_243528# a_403521_244568# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X35 a_395162_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X36 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X37 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X38 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X39 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X40 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X41 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X42 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X43 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X44 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X45 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X46 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X47 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X48 a_402731_244568# a_401151_244568# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X49 a_365708_259299# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X50 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X51 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X52 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X53 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X54 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X55 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X56 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X57 a_409498_256643# a_404041_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X58 a_395682_259299# a_383940_262205# a_395162_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X59 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X60 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X61 a_409618_260539# a_404041_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X62 a_401941_244568# a_401151_244568# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X63 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X64 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X65 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X66 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X67 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X68 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X69 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X70 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X71 a_409618_260539# a_404041_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X72 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X73 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X74 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X75 a_411044_242557# a_402461_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X76 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X77 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X78 a_401151_244568# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X79 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X80 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X81 a_402461_244568# a_402461_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X82 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X83 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X84 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X85 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X86 a_404041_244568# a_409618_256263# a_409618_260539# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X87 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X88 a_404831_244568# a_401271_243528# a_404311_244568# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X89 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X90 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X91 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X92 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X93 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X94 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X95 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X96 a_401271_243528# a_401271_243528# a_401151_244568# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X97 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X98 a_403521_244568# a_401151_244568# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X99 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X100 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X101 a_410724_251737# a_410134_251737# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X102 a_409618_256263# a_409498_256643# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X103 a_411044_251737# a_403251_244568# a_410724_251737# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X104 a_409818_256643# a_409618_256263# a_409498_256643# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X105 a_386992_259299# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X106 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X107 a_410134_251737# a_410134_251737# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X108 a_403251_244568# a_403251_244568# a_410134_251737# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X109 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X110 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X111 a_409818_256643# a_409618_256263# a_409498_256643# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X112 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X113 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X114 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X115 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X116 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X117 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X118 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X119 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X120 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X121 a_383620_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X122 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X123 a_373878_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X124 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X125 a_409498_256643# a_404041_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X126 a_401151_244568# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X127 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X128 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X129 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X130 a_403251_244568# a_401271_243528# a_402731_244568# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X131 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X132 a_383940_262205# a_374398_259299# a_383620_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X133 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
C0 a_401941_244568# a_404831_244568# 0.13684f
C1 a_403521_244568# a_402731_244568# 0.84407f
C2 a_409618_256263# a_404041_244568# 1.45171f
C3 a_404041_244568# a_403251_244568# 0.33183f
C4 a_365828_265695# a_365708_259299# 0.74385f
C5 a_404041_244568# a_409618_260539# 3.00275f
C6 a_403521_244568# a_401941_244568# 0.34178f
C7 a_365828_265695# a_402731_244568# 0.0069f
C8 a_401941_244568# a_365828_265695# 0.00563f
C9 a_404041_244568# w_364522_258756# 1.72336f
C10 a_365828_265695# a_365828_259091# 0.00331f
C11 a_373878_259299# a_365708_259299# 0.98664f
C12 a_404311_244568# a_402731_244568# 0.30154f
C13 a_404311_244568# a_401941_244568# 0.30103f
C14 a_373878_259299# a_365828_259091# 0.99903f
C15 a_386992_259299# a_365828_265695# 0.7554f
C16 a_410724_251737# a_411044_251737# 1.15251f
C17 a_410134_251737# a_411044_251737# 0.0849f
C18 a_401271_243528# a_402731_244568# 0.63243f
C19 a_410134_251737# a_410724_251737# 0.36588f
C20 a_411044_242557# a_402461_244568# 0.20751f
C21 a_401941_244568# a_401271_243528# 2.86501f
C22 a_404041_244568# a_404831_244568# 2.48301f
C23 a_374398_259299# a_365708_259299# 0.07017f
C24 a_404041_244568# a_403521_244568# 2.39829f
C25 a_411044_251737# a_403251_244568# 0.2042f
C26 a_365828_259091# a_374398_259299# 0.50349f
C27 a_410724_251737# a_403251_244568# 1.45997f
C28 a_409498_256643# a_409818_256643# 2.17202f
C29 a_410134_251737# a_403251_244568# 1.85176f
C30 a_401151_244568# a_402461_244568# 0.13364f
C31 w_364522_258756# a_383940_262205# 15.504f
C32 a_409618_256263# a_409818_256643# 0.57687f
C33 a_409818_256643# a_409618_260539# 0.0136f
C34 a_404311_244568# a_404041_244568# 2.29591f
C35 a_401151_244568# a_403251_244568# 0.13521f
C36 a_409618_256263# a_409498_256643# 3.29507f
C37 a_409498_256643# a_409618_260539# 0.36393f
C38 a_395682_259299# a_383940_262205# 0.50349f
C39 a_403251_244568# a_402461_244568# 0.58599f
C40 a_401151_244568# w_364522_258756# 44.8668f
C41 a_386992_259299# a_395162_259299# 0.98664f
C42 a_401941_244568# a_402731_244568# 0.84535f
C43 a_409618_256263# a_409618_260539# 3.58908f
C44 a_365828_259091# a_365708_259299# 29.489f
C45 w_364522_258756# a_402461_244568# 1.21291f
C46 a_403251_244568# w_364522_258756# 1.12778f
C47 a_404041_244568# a_401271_243528# 0.62193f
C48 a_383620_262205# a_383940_262205# 1.13981f
C49 a_395682_259299# w_364522_258756# 1.49117f
C50 a_365828_265695# a_383940_262205# 0.01792f
C51 a_401151_244568# a_404831_244568# 0.98673f
C52 a_401151_244568# a_403521_244568# 1.46461f
C53 a_404831_244568# a_402461_244568# 0.08091f
C54 a_401151_244568# a_365828_265695# 2.15734f
C55 a_409618_256263# a_404831_244568# 0.12451f
C56 a_403521_244568# a_402461_244568# 0.10043f
C57 a_404041_244568# a_402731_244568# 0.17025f
C58 a_403251_244568# a_404831_244568# 0.08038f
C59 a_404831_244568# a_409618_260539# 0
C60 a_403251_244568# a_403521_244568# 2.29847f
C61 a_404041_244568# a_401941_244568# 0.17047f
C62 w_364522_258756# a_404831_244568# 2.87066f
C63 a_403521_244568# w_364522_258756# 7.51371f
C64 a_401151_244568# a_404311_244568# 2.37681f
C65 w_364522_258756# a_365828_265695# 19.3145f
C66 a_404311_244568# a_402461_244568# 0.10003f
C67 a_383620_262205# a_377450_262205# 0.52252f
C68 a_404311_244568# a_403251_244568# 0.10042f
C69 a_374398_259299# a_383940_262205# 0.28491f
C70 a_373878_259299# w_364522_258756# 3.05677f
C71 a_404311_244568# w_364522_258756# 6.35462f
C72 a_401151_244568# a_401271_243528# 3.41485f
C73 a_383940_262205# a_395162_259299# 0.99903f
C74 a_401271_243528# a_402461_244568# 0.63416f
C75 a_403251_244568# a_401271_243528# 0.62309f
C76 a_403521_244568# a_404831_244568# 0.13662f
C77 w_364522_258756# a_401271_243528# 14.5258f
C78 a_403521_244568# a_365828_265695# 0.00915f
C79 w_364522_258756# a_374398_259299# 1.76606f
C80 w_364522_258756# a_395162_259299# 3.05677f
C81 a_401151_244568# a_402731_244568# 1.46427f
C82 a_404311_244568# a_404831_244568# 2.35844f
C83 a_401151_244568# a_401941_244568# 1.80913f
C84 a_404311_244568# a_403521_244568# 0.80509f
C85 a_402731_244568# a_402461_244568# 2.30103f
C86 a_395682_259299# a_395162_259299# 0.8533f
C87 a_373878_259299# a_365828_265695# 0
C88 a_404311_244568# a_365828_265695# 0.28741f
C89 a_401941_244568# a_402461_244568# 2.41261f
C90 a_403251_244568# a_402731_244568# 2.40482f
C91 a_386992_259299# a_383940_262205# 29.4825f
C92 a_403251_244568# a_401941_244568# 0.17152f
C93 w_364522_258756# a_365708_259299# 48.8544f
C94 a_377450_262205# a_374398_259299# 36.6185f
C95 w_364522_258756# a_402731_244568# 7.43186f
C96 a_401271_243528# a_404831_244568# 0.54995f
C97 a_383620_262205# a_374398_259299# 0.86502f
C98 a_401941_244568# w_364522_258756# 7.43338f
C99 a_403521_244568# a_401271_243528# 0.62333f
C100 w_364522_258756# a_365828_259091# 16.3092f
C101 a_365828_265695# a_374398_259299# 0.01878f
C102 a_365828_265695# a_395162_259299# 0
C103 a_386992_259299# w_364522_258756# 48.8285f
C104 a_404311_244568# a_401271_243528# 0.62105f
C105 a_409818_256643# a_404041_244568# 0.00933f
C106 a_401151_244568# a_404041_244568# 0.59986f
C107 a_409498_256643# a_404041_244568# 0.85546f
C108 a_373878_259299# a_374398_259299# 0.91714f
C109 a_395682_259299# a_386992_259299# 0.06695f
C110 a_404831_244568# a_402731_244568# 0.13558f
C111 a_404041_244568# a_402461_244568# 0.10021f
C112 a_411044_242557# a_376520_259212# 6.1069f
C113 a_411044_251737# a_376520_259212# 4.75873f
C114 a_410724_251737# a_376520_259212# 2.90137f
C115 a_410134_251737# a_376520_259212# 6.39712f
C116 a_409818_256643# a_376520_259212# 5.97383f
C117 a_409498_256643# a_376520_259212# 8.54632f
C118 a_409618_256263# a_376520_259212# 12.5882f
C119 a_409618_260539# a_376520_259212# 7.6582f
C120 a_404831_244568# a_376520_259212# 10.5405f
C121 a_404041_244568# a_376520_259212# 11.5785f
C122 a_403251_244568# a_376520_259212# 5.05938f
C123 a_402461_244568# a_376520_259212# 7.97268f
C124 a_401271_243528# a_376520_259212# 2.45016f
C125 a_404311_244568# a_376520_259212# 0.15844f
C126 a_403521_244568# a_376520_259212# 0.03326f
C127 a_402731_244568# a_376520_259212# 0.03284f
C128 a_401941_244568# a_376520_259212# 0.03295f
C129 a_401151_244568# a_376520_259212# 2.60775f
C130 a_395682_259299# a_376520_259212# 0.40915f
C131 a_395162_259299# a_376520_259212# 0.29295f
C132 a_383940_262205# a_376520_259212# 4.92556f
C133 a_383620_262205# a_376520_259212# 2.7563f
C134 a_377450_262205# a_376520_259212# 40.1477f
C135 a_374398_259299# a_376520_259212# 12.9247f
C136 a_365828_259091# a_376520_259212# 25.3712f
C137 a_373878_259299# a_376520_259212# 0.20081f
C138 a_386992_259299# a_376520_259212# 3.24772f
C139 a_365708_259299# a_376520_259212# 3.20723f
C140 a_365828_265695# a_376520_259212# 24.117f
C141 w_364522_258756# a_376520_259212# 0.94999p
.ends

.subckt TOP CCM_OUT PU VDD VSS VIN_OUT BCM_OUT VCM_OUT VIN VBIAS EN PD
Xsc_tieh_tiel$1_0 PD PU sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157#
+ VDD sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# VSS sc_tieh_tiel$1
Xio_secondary_5p0$1_0 EN m3_419992_265695# VSS VDD io_secondary_5p0$1
XM_0 M_0/a_402461_244568# M_0/a_410134_251737# VSS M_0/a_403521_244568# a_499016_248165#
+ BCM_OUT m4_400150_261569# M_0/a_409618_260539# VIN_OUT a_498947_268180# CCM_OUT
+ M_0/a_403251_244568# m3_419992_265695# M_0/a_404311_244568# VSS M_0/a_401941_244568#
+ m4_400150_261569# M_0/a_404041_244568# M_0/a_409498_256643# M_0/a_402731_244568#
+ M_0/a_401151_244568# VCM_OUT VDD M
D0 a_498947_268180# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D1 a_498947_268180# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D2 VSS a_499016_248165# diode_nd2ps_06v0 pj=40u area=99.99999p
X0 a_498947_268180# VIN VDD ppolyf_u r_width=40u r_length=10u
D3 a_499016_248165# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D4 a_499016_248165# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D5 VSS a_499016_248165# diode_nd2ps_06v0 pj=40u area=99.99999p
D6 a_498947_268180# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D7 VSS a_498947_268180# diode_nd2ps_06v0 pj=40u area=99.99999p
D8 a_499016_248165# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D9 a_499016_248165# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D10 VSS a_498947_268180# diode_nd2ps_06v0 pj=40u area=99.99999p
D11 VSS a_499016_248165# diode_nd2ps_06v0 pj=40u area=99.99999p
D12 VSS a_498947_268180# diode_nd2ps_06v0 pj=40u area=99.99999p
D13 a_498947_268180# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
X1 a_499016_248165# VBIAS VDD ppolyf_u r_width=40u r_length=10u
D14 VSS a_499016_248165# diode_nd2ps_06v0 pj=40u area=99.99999p
D15 VSS a_498947_268180# diode_nd2ps_06v0 pj=40u area=99.99999p
C0 TEXT$22_0/m2_7200_0# TEXT$9_0/m1_2880_0# 0
C1 TEXT$1_0/m1_6000_0# TEXT$1_0/m1_7200_0# 0.2838f
C2 TEXT$21_0/m4_10800_0# TEXT$21_0/m4_11700_0# 0.14096f
C3 TEXT$24_0/m3_960_0# TEXT$9_0/m1_2160_0# 0
C4 TEXT$24_0/m3_2160_0# TEXT$9_0/m1_960_0# 0
C5 sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# PD 0.00624f
C6 TEXT$21_0/m4_2160_0# TEXT$22_0/m2_1440_0# 0
C7 TEXT$1_0/m1_2400_0# TEXT$6_0/m4_2400_0# 0.00679f
C8 TEXT$3_0/m2_4800_0# TEXT$20_0/m3_7920_720# 0
C9 TEXT$24_0/m3_9600_0# TEXT$9_0/m1_9600_0# 0.01567f
C10 TEXT$24_0/m3_5760_0# TEXT$21_0/m4_9360_0# 0
C11 TEXT$21_0/m4_7920_720# TEXT$9_0/m1_3840_0# -0
C12 M_0/a_409618_260539# m4_400150_261569# -0
C13 TEXT$24_0/m3_5760_0# TEXT$7_0/m2_4800_960# 0.00343f
C14 TEXT$23_0/m1_1440_0# TEXT$22_0/m2_720_0# 0.00168f
C15 TEXT$20_0/m3_7200_0# TEXT$20_0/m3_7920_720# 0.12093f
C16 TEXT$8_0/m4_6720_0# TEXT$20_0/m3_10800_0# 0
C17 TEXT$23_0/m1_3780_0# TEXT$20_0/m3_3780_0# 0.00157f
C18 TEXT$22_0/m2_9360_0# TEXT$20_0/m3_9360_0# 0.42195f
C19 TEXT$21_0/m4_16560_0# TEXT$21_0/m4_17280_0# 0.15155f
C20 TEXT$24_0/m3_10560_0# TEXT$20_0/m3_14400_0# 0.01775f
C21 TEXT$23_0/m1_5760_0# TEXT$1_0/m1_3600_0# 0.00988f
C22 TEXT$21_0/m4_10080_0# TEXT$20_0/m3_10080_0# 0.40607f
C23 TEXT$22_0/m2_5760_0# TEXT$6_0/m4_3600_0# 0
C24 TEXT$23_0/m1_7920_720# TEXT$23_0/m1_7200_0# 0.10344f
C25 TEXT$23_0/m1_10800_0# TEXT$20_0/m3_10800_0# 0.0029f
C26 TEXT$8_0/m4_10560_0# TEXT$9_0/m1_9600_0# -0
C27 TEXT$24_0/m3_3840_0# TEXT$22_0/m2_8640_0# 0.00169f
C28 TEXT$4_0/m3_7200_0# TEXT$22_0/m2_9360_0# 0
C29 TEXT$21_0/m4_1440_0# TEXT$20_0/m3_1440_0# 0.36769f
C30 TEXT$23_0/m1_6480_0# TEXT$6_0/m4_3600_0# 0
C31 TEXT$3_0/m2_0_0# TEXT$23_0/m1_2880_720# 0
C32 TEXT$4_0/m3_7200_0# TEXT$1_0/m1_6000_0# 0.00242f
C33 TEXT$24_0/m3_4800_960# TEXT$21_0/m4_9360_0# 0
C34 TEXT$24_0/m3_9600_0# TEXT$23_0/m1_13680_0# 0
C35 TEXT$24_0/m3_4800_960# TEXT$7_0/m2_4800_960# 0.42246f
C36 TEXT$21_0/m4_16560_0# TEXT$20_0/m3_16560_0# 0.40081f
C37 TEXT$23_0/m1_14400_0# TEXT$9_0/m1_10560_0# 0.01107f
C38 TEXT$4_0/m3_0_0# TEXT$21_0/m4_2160_0# 0
C39 TEXT$22_0/m2_9360_0# TEXT$3_0/m2_7200_0# 0.01999f
C40 TEXT$23_0/m1_2880_720# TEXT$20_0/m3_3780_0# 0
C41 TEXT$23_0/m1_3780_0# TEXT$20_0/m3_2880_720# 0
C42 TEXT$9_0/m1_5760_0# TEXT$8_0/m4_5760_0# 0.00251f
C43 TEXT$8_0/m4_10560_0# TEXT$20_0/m3_15120_0# 0
C44 TEXT$1_0/m1_10800_0# TEXT$3_0/m2_10800_0# 1.16108f
C45 TEXT$7_0/m2_9600_0# TEXT$7_0/m2_10560_0# 0.13915f
C46 TEXT$20_0/m3_12960_0# TEXT$3_0/m2_10800_0# 0
C47 TEXT$1_0/m1_6000_0# TEXT$3_0/m2_7200_0# 0.007f
C48 TEXT$22_0/m2_17280_0# TEXT$22_0/m2_18000_0# 0.17402f
C49 TEXT$9_0/m1_4800_960# TEXT$7_0/m2_5760_0# 0
C50 TEXT$3_0/m2_2400_0# TEXT$6_0/m4_2400_0# 0.00713f
C51 TEXT$20_0/m3_8640_0# TEXT$20_0/m3_9360_0# 0.26159f
C52 TEXT$8_0/m4_960_0# TEXT$24_0/m3_0_0# 0
C53 TEXT$9_0/m1_960_0# TEXT$9_0/m1_2160_0# 0.1022f
C54 TEXT$21_0/m4_15840_0# TEXT$23_0/m1_15840_0# 0
C55 TEXT$23_0/m1_10080_0# TEXT$23_0/m1_9360_0# 0.1367f
C56 TEXT$23_0/m1_15120_0# TEXT$20_0/m3_15120_0# 0.0029f
C57 VIN_OUT m4_400150_261569# 0.03198f
C58 TEXT$9_0/m1_6720_0# TEXT$7_0/m2_5760_0# 0.00386f
C59 TEXT$22_0/m2_13680_0# TEXT$9_0/m1_9600_0# 0
C60 TEXT$23_0/m1_1440_0# TEXT$22_0/m2_1440_0# 0.36465f
C61 TEXT$23_0/m1_720_0# TEXT$20_0/m3_720_0# 0.00233f
C62 TEXT$24_0/m3_3840_0# TEXT$22_0/m2_7920_720# 0
C63 TEXT$8_0/m4_5760_0# TEXT$8_0/m4_6720_0# 0.22111f
C64 TEXT$8_0/m4_2880_0# TEXT$20_0/m3_7200_0# 0.00108f
C65 TEXT$24_0/m3_2880_0# TEXT$24_0/m3_2160_0# 0.14271f
C66 TEXT$23_0/m1_11700_0# TEXT$3_0/m2_9600_0# 0
C67 TEXT$22_0/m2_8640_0# TEXT$9_0/m1_3840_0# 0.00207f
C68 TEXT$23_0/m1_5760_0# TEXT$3_0/m2_3600_0# 0
C69 TEXT$24_0/m3_7680_0# VDD 0.00386f
C70 TEXT$4_0/m3_6000_0# TEXT$4_0/m3_7200_0# 0.31804f
C71 TEXT$8_0/m4_6720_0# TEXT$7_0/m2_6720_0# 0.01464f
C72 TEXT$23_0/m1_2880_720# TEXT$20_0/m3_2880_720# 0.00212f
C73 TEXT$22_0/m2_15120_0# TEXT$21_0/m4_15120_0# 0.00342f
C74 TEXT$22_0/m2_9360_0# TEXT$8_0/m4_4800_960# 0
C75 TEXT$7_0/m2_7680_0# TEXT$20_0/m3_11700_0# 0
C76 TEXT$9_0/m1_10560_0# VDD 0.03368f
C77 TEXT$22_0/m2_15120_0# TEXT$1_0/m1_12000_0# 0
C78 TEXT$21_0/m4_9360_0# TEXT$9_0/m1_4800_960# 0
C79 TEXT$22_0/m2_14400_0# TEXT$20_0/m3_14400_0# 0.41009f
C80 TEXT$9_0/m1_4800_960# TEXT$7_0/m2_4800_960# 0.42103f
C81 TEXT$8_0/m4_3840_0# TEXT$8_0/m4_4800_960# 0.15822f
C82 TEXT$4_0/m3_10800_0# TEXT$3_0/m2_10800_0# 1.15603f
C83 TEXT$6_0/m4_9600_0# TEXT$3_0/m2_10800_0# 0
C84 TEXT$6_0/m4_10800_0# TEXT$3_0/m2_9600_0# 0
C85 TEXT$21_0/m4_10080_0# TEXT$9_0/m1_5760_0# 0
C86 TEXT$22_0/m2_10080_0# TEXT$22_0/m2_10800_0# 0.20701f
C87 TEXT$23_0/m1_2160_0# TEXT$22_0/m2_1440_0# 0
C88 TEXT$23_0/m1_10800_0# TEXT$7_0/m2_6720_0# 0
C89 TEXT$21_0/m4_14400_0# TEXT$8_0/m4_9600_0# 0.01f
C90 sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# VDD 0.00261f
C91 TEXT$21_0/m4_2160_0# TEXT$23_0/m1_1440_0# 0
C92 TEXT$22_0/m2_13680_0# TEXT$23_0/m1_13680_0# 0.34645f
C93 TEXT$21_0/m4_11700_0# TEXT$22_0/m2_10800_0# 0
C94 TEXT$3_0/m2_6000_0# TEXT$3_0/m2_7200_0# 0.25104f
C95 TEXT$22_0/m2_7920_720# TEXT$9_0/m1_3840_0# 0
C96 TEXT$21_0/m4_11700_0# TEXT$1_0/m1_8400_0# 0
C97 TEXT$1_0/m1_7200_0# TEXT$1_0/m1_8400_0# 0.09175f
C98 TEXT$21_0/m4_11700_0# TEXT$21_0/m4_12960_0# 0.02736f
C99 TEXT$24_0/m3_2160_0# TEXT$9_0/m1_2880_0# 0
C100 TEXT$24_0/m3_5760_0# TEXT$22_0/m2_9360_0# 0
C101 TEXT$22_0/m2_2160_0# TEXT$20_0/m3_1440_0# 0
C102 TEXT$22_0/m2_1440_0# TEXT$20_0/m3_2160_0# 0.00148f
C103 TEXT$21_0/m4_10800_0# TEXT$20_0/m3_11700_0# 0
C104 TEXT$1_0/m1_3600_0# TEXT$6_0/m4_3600_0# 0.0042f
C105 TEXT$21_0/m4_2880_720# TEXT$22_0/m2_2160_0# 0
C106 TEXT$21_0/m4_2880_720# TEXT$21_0/m4_3780_0# 0.10067f
C107 TEXT$8_0/m4_4800_960# TEXT$20_0/m3_8640_0# 0
C108 TEXT$24_0/m3_10560_0# TEXT$9_0/m1_10560_0# 0.01345f
C109 TEXT$4_0/m3_0_0# TEXT$22_0/m2_2880_720# 0
C110 TEXT$22_0/m2_15120_0# TEXT$4_0/m3_12000_0# 0
C111 TEXT$22_0/m2_14400_0# TEXT$6_0/m4_12000_0# 0
C112 TEXT$4_0/m3_1200_0# TEXT$21_0/m4_3780_0# 0
C113 TEXT$24_0/m3_2880_0# TEXT$9_0/m1_2160_0# 0
C114 TEXT$21_0/m4_10080_0# TEXT$23_0/m1_10800_0# -0
C115 TEXT$22_0/m2_2160_0# TEXT$1_0/m1_0_0# 0
C116 TEXT$21_0/m4_8640_0# TEXT$23_0/m1_8640_0# 0
C117 TEXT$23_0/m1_1440_0# TEXT$23_0/m1_720_0# 0.30936f
C118 TEXT$22_0/m2_10080_0# TEXT$20_0/m3_10080_0# 0.40884f
C119 TEXT$21_0/m4_17280_0# TEXT$20_0/m3_16560_0# 0
C120 TEXT$23_0/m1_8640_0# TEXT$7_0/m2_3840_0# 0
C121 TEXT$21_0/m4_2160_0# TEXT$23_0/m1_2160_0# -0
C122 TEXT$1_0/m1_7200_0# TEXT$20_0/m3_10080_0# 0
C123 TEXT$8_0/m4_10560_0# TEXT$24_0/m3_9600_0# 0.00253f
C124 TEXT$4_0/m3_0_0# TEXT$23_0/m1_2160_0# 0
C125 TEXT$23_0/m1_4320_0# TEXT$22_0/m2_3780_0# 0
C126 TEXT$24_0/m3_4800_960# TEXT$22_0/m2_9360_0# 0
C127 TEXT$21_0/m4_7920_720# TEXT$6_0/m4_4800_0# 0.01309f
C128 VDD EN 2.4043f
C129 TEXT$21_0/m4_2160_0# TEXT$20_0/m3_2160_0# 0.4f
C130 TEXT$4_0/m3_8400_0# TEXT$21_0/m4_11700_0# 0
C131 TEXT$4_0/m3_8400_0# TEXT$1_0/m1_7200_0# 0
C132 TEXT$24_0/m3_4800_960# TEXT$8_0/m4_3840_0# 0.00215f
C133 TEXT$24_0/m3_10560_0# TEXT$23_0/m1_14400_0# 0
C134 TEXT$21_0/m4_10800_0# TEXT$6_0/m4_8400_0# 0.03468f
C135 TEXT$4_0/m3_3600_0# TEXT$6_0/m4_3600_0# 1.10156f
C136 TEXT$4_0/m3_0_0# TEXT$20_0/m3_2160_0# 0.0125f
C137 TEXT$22_0/m2_2880_720# TEXT$22_0/m2_3780_0# 0.06867f
C138 TEXT$24_0/m3_2880_0# TEXT$8_0/m4_2880_0# 0.66142f
C139 TEXT$21_0/m4_4320_0# TEXT$22_0/m2_3780_0# 0
C140 TEXT$24_0/m3_2160_0# TEXT$23_0/m1_5760_0# 0
C141 TEXT$21_0/m4_15120_0# TEXT$3_0/m2_12000_0# 0
C142 TEXT$1_0/m1_12000_0# TEXT$3_0/m2_12000_0# 1.12229f
C143 TEXT$21_0/m4_11700_0# TEXT$3_0/m2_8400_0# 0
C144 TEXT$1_0/m1_7200_0# TEXT$3_0/m2_8400_0# 0.00181f
C145 TEXT$3_0/m2_3600_0# TEXT$6_0/m4_3600_0# 0.00883f
C146 TEXT$20_0/m3_9360_0# TEXT$20_0/m3_10080_0# 0.12171f
C147 TEXT$8_0/m4_960_0# TEXT$24_0/m3_2160_0# 0.00171f
C148 TEXT$9_0/m1_2160_0# TEXT$9_0/m1_2880_0# 0.1022f
C149 TEXT$21_0/m4_16560_0# TEXT$23_0/m1_16560_0# -0
C150 TEXT$4_0/m3_1200_0# TEXT$1_0/m1_0_0# 0.00156f
C151 TEXT$24_0/m3_6720_0# TEXT$7_0/m2_5760_0# 0.00701f
C152 TEXT$22_0/m2_13680_0# TEXT$24_0/m3_9600_0# 0
C153 TEXT$6_0/m4_3600_0# TEXT$20_0/m3_6480_0# 0
C154 TEXT$23_0/m1_15840_0# TEXT$20_0/m3_15840_0# 0.00322f
C155 TEXT$9_0/m1_7680_0# TEXT$7_0/m2_6720_0# 0.00567f
C156 TEXT$22_0/m2_14400_0# TEXT$9_0/m1_10560_0# 0
C157 TEXT$8_0/m4_10560_0# TEXT$23_0/m1_15120_0# 0
C158 TEXT$21_0/m4_4320_0# TEXT$23_0/m1_4320_0# -0.00759f
C159 TEXT$4_0/m3_7200_0# TEXT$20_0/m3_10080_0# 0.019f
C160 TEXT$24_0/m3_4800_960# TEXT$20_0/m3_8640_0# 0.01605f
C161 TEXT$22_0/m2_2160_0# TEXT$3_0/m2_0_0# 0.00873f
C162 TEXT$23_0/m1_12960_0# TEXT$3_0/m2_10800_0# 0
C163 TEXT$22_0/m2_9360_0# TEXT$9_0/m1_4800_960# 0
C164 TEXT$24_0/m3_10560_0# VDD 0.00927f
C165 TEXT$4_0/m3_7200_0# TEXT$4_0/m3_8400_0# 0.12422f
C166 TEXT$21_0/m4_14400_0# TEXT$7_0/m2_9600_0# 0
C167 TEXT$21_0/m4_3780_0# TEXT$20_0/m3_3780_0# 0.19343f
C168 TEXT$3_0/m2_7200_0# TEXT$20_0/m3_10080_0# 0
C169 TEXT$22_0/m2_15840_0# TEXT$21_0/m4_15840_0# 0.00404f
C170 TEXT$24_0/m3_2880_0# TEXT$24_0/m3_3840_0# 0.14642f
C171 TEXT$9_0/m1_7680_0# TEXT$8_0/m4_9600_0# 0
C172 TEXT$22_0/m2_15120_0# TEXT$20_0/m3_15120_0# 0.36742f
C173 TEXT$9_0/m1_4800_960# TEXT$8_0/m4_3840_0# -0
C174 TEXT$7_0/m2_2880_0# TEXT$23_0/m1_7200_0# 0
C175 TEXT$23_0/m1_2160_0# TEXT$23_0/m1_1440_0# 0.13524f
C176 TEXT$22_0/m2_10080_0# TEXT$9_0/m1_5760_0# 0
C177 TEXT$4_0/m3_1200_0# TEXT$22_0/m2_4320_0# 0
C178 TEXT$9_0/m1_2880_0# TEXT$8_0/m4_2880_0# 0.00298f
C179 TEXT$8_0/m4_7680_0# TEXT$8_0/m4_6720_0# 0.30955f
C180 TEXT$22_0/m2_11700_0# TEXT$3_0/m2_9600_0# 0.00166f
C181 TEXT$4_0/m3_12000_0# TEXT$3_0/m2_12000_0# 1.1133f
C182 TEXT$4_0/m3_7200_0# TEXT$3_0/m2_8400_0# 0
C183 TEXT$6_0/m4_12000_0# TEXT$3_0/m2_10800_0# 0
C184 TEXT$6_0/m4_10800_0# TEXT$3_0/m2_12000_0# 0
C185 TEXT$21_0/m4_10800_0# TEXT$9_0/m1_6720_0# 0
C186 TEXT$22_0/m2_3780_0# TEXT$1_0/m1_1200_0# 0
C187 TEXT$23_0/m1_11700_0# TEXT$7_0/m2_7680_0# 0
C188 TEXT$8_0/m4_9600_0# TEXT$20_0/m3_14400_0# 0
C189 TEXT$22_0/m2_14400_0# TEXT$23_0/m1_14400_0# 0.40648f
C190 TEXT$7_0/m2_0_0# VDD 0.02935f
C191 TEXT$22_0/m2_10800_0# TEXT$20_0/m3_11700_0# 0
C192 TEXT$3_0/m2_7200_0# TEXT$3_0/m2_8400_0# 0.0908f
C193 TEXT$21_0/m4_2880_720# TEXT$3_0/m2_0_0# 0
C194 TEXT$4_0/m3_2400_0# TEXT$23_0/m1_4320_0# 0
C195 TEXT$21_0/m4_11700_0# TEXT$8_0/m4_6720_0# 0.00103f
C196 TEXT$1_0/m1_8400_0# TEXT$1_0/m1_9600_0# 0.27287f
C197 TEXT$21_0/m4_12960_0# TEXT$21_0/m4_13680_0# 0.20695f
C198 TEXT$9_0/m1_4800_960# TEXT$20_0/m3_8640_0# 0
C199 TEXT$21_0/m4_11700_0# TEXT$20_0/m3_12960_0# 0
C200 TEXT$22_0/m2_2160_0# TEXT$20_0/m3_2880_720# 0.00104f
C201 TEXT$1_0/m1_8400_0# TEXT$20_0/m3_11700_0# 0
C202 TEXT$21_0/m4_12960_0# TEXT$20_0/m3_11700_0# 0
C203 TEXT$1_0/m1_4800_0# TEXT$6_0/m4_4800_0# 0.00618f
C204 TEXT$8_0/m4_960_0# TEXT$9_0/m1_2160_0# 0
C205 TEXT$23_0/m1_4320_0# TEXT$1_0/m1_1200_0# 0.00758f
C206 TEXT$21_0/m4_2880_720# TEXT$20_0/m3_3780_0# 0
C207 TEXT$21_0/m4_3780_0# TEXT$20_0/m3_2880_720# 0
C208 TEXT$21_0/m4_7200_0# TEXT$23_0/m1_7200_0# 0
C209 TEXT$6_0/m4_0_0# TEXT$6_0/m4_1200_0# 0.26602f
C210 TEXT$23_0/m1_6480_0# TEXT$23_0/m1_7200_0# 0.29377f
C211 TEXT$1_0/m1_0_0# TEXT$3_0/m2_0_0# 1.13089f
C212 TEXT$4_0/m3_1200_0# TEXT$20_0/m3_3780_0# 0.0104f
C213 TEXT$4_0/m3_2400_0# TEXT$21_0/m4_4320_0# 0
C214 TEXT$22_0/m2_8640_0# TEXT$23_0/m1_8640_0# 0.40245f
C215 TEXT$22_0/m2_10080_0# TEXT$23_0/m1_10800_0# 0.00198f
C216 TEXT$24_0/m3_3840_0# TEXT$9_0/m1_2880_0# 0.00155f
C217 TEXT$21_0/m4_11700_0# TEXT$23_0/m1_10800_0# 0
C218 TEXT$24_0/m3_3840_0# TEXT$8_0/m4_4800_960# 0
C219 TEXT$21_0/m4_4320_0# TEXT$1_0/m1_1200_0# 0
C220 TEXT$21_0/m4_17280_0# TEXT$20_0/m3_18000_0# 0
C221 TEXT$23_0/m1_2160_0# TEXT$20_0/m3_2160_0# 0.00218f
C222 TEXT$22_0/m2_7920_720# TEXT$6_0/m4_4800_0# 0
C223 TEXT$23_0/m1_4320_0# TEXT$22_0/m2_5760_0# 0
C224 TEXT$22_0/m2_4320_0# TEXT$7_0/m2_0_0# 0.01201f
C225 TEXT$24_0/m3_5760_0# TEXT$20_0/m3_10080_0# 0.02608f
C226 TEXT$22_0/m2_10800_0# TEXT$6_0/m4_8400_0# 0
C227 TEXT$22_0/m2_3780_0# TEXT$3_0/m2_1200_0# 0.00714f
C228 TEXT$21_0/m4_2880_720# TEXT$20_0/m3_2880_720# 0.23623f
C229 TEXT$4_0/m3_8400_0# TEXT$1_0/m1_9600_0# 0
C230 TEXT$21_0/m4_17280_0# TEXT$23_0/m1_16560_0# 0
C231 TEXT$4_0/m3_9600_0# TEXT$1_0/m1_8400_0# 0.00258f
C232 TEXT$23_0/m1_7920_720# TEXT$22_0/m2_7200_0# 0
C233 TEXT$4_0/m3_8400_0# TEXT$20_0/m3_11700_0# 0
C234 TEXT$21_0/m4_11700_0# TEXT$6_0/m4_9600_0# 0.00175f
C235 TEXT$4_0/m3_4800_0# TEXT$6_0/m4_4800_0# 1.10696f
C236 TEXT$1_0/m1_8400_0# TEXT$6_0/m4_8400_0# 0.00466f
C237 TEXT$8_0/m4_0_0# TEXT$23_0/m1_4320_0# -0
C238 TEXT$22_0/m2_7920_720# TEXT$23_0/m1_8640_0# 0
C239 TEXT$22_0/m2_4320_0# TEXT$20_0/m3_3780_0# 0
C240 TEXT$22_0/m2_3780_0# TEXT$20_0/m3_4320_0# 0
C241 TEXT$21_0/m4_4320_0# TEXT$22_0/m2_5760_0# 0
C242 TEXT$21_0/m4_5760_0# TEXT$22_0/m2_4320_0# 0
C243 TEXT$21_0/m4_9360_0# TEXT$23_0/m1_9360_0# -0
C244 TEXT$23_0/m1_9360_0# TEXT$7_0/m2_4800_960# 0
C245 TEXT$23_0/m1_10080_0# TEXT$7_0/m2_5760_0# 0.00141f
C246 TEXT$1_0/m1_0_0# TEXT$20_0/m3_2880_720# 0
C247 TEXT$1_0/m1_9600_0# TEXT$3_0/m2_8400_0# 0
C248 TEXT$20_0/m3_15120_0# TEXT$3_0/m2_12000_0# 0
C249 TEXT$21_0/m4_5760_0# TEXT$21_0/m4_6480_0# 0.18409f
C250 TEXT$3_0/m2_8400_0# TEXT$20_0/m3_11700_0# 0
C251 TEXT$3_0/m2_4800_0# TEXT$6_0/m4_4800_0# 0.00754f
C252 TEXT$23_0/m1_4320_0# TEXT$3_0/m2_1200_0# 0
C253 TEXT$9_0/m1_2880_0# TEXT$9_0/m1_3840_0# 0.13265f
C254 VDD TEXT$7_0/m2_3840_0# 0.03406f
C255 TEXT$4_0/m3_2400_0# TEXT$1_0/m1_1200_0# 0.00242f
C256 TEXT$8_0/m4_0_0# TEXT$21_0/m4_4320_0# 0.01821f
C257 TEXT$9_0/m1_3840_0# TEXT$8_0/m4_4800_960# 0
C258 TEXT$24_0/m3_7680_0# TEXT$7_0/m2_6720_0# 0.01136f
C259 TEXT$22_0/m2_14400_0# TEXT$24_0/m3_10560_0# 0
C260 TEXT$23_0/m1_16560_0# TEXT$20_0/m3_16560_0# 0.00203f
C261 TEXT$9_0/m1_7680_0# TEXT$7_0/m2_9600_0# 0
C262 TEXT$9_0/m1_9600_0# TEXT$7_0/m2_7680_0# 0
C263 TEXT$23_0/m1_4320_0# TEXT$20_0/m3_4320_0# 0.00213f
C264 TEXT$9_0/m1_5760_0# TEXT$8_0/m4_4800_960# 0
C265 TEXT$9_0/m1_7680_0# TEXT$8_0/m4_7680_0# 0
C266 TEXT$21_0/m4_4320_0# TEXT$3_0/m2_1200_0# 0
C267 VDD TEXT$8_0/m4_2160_0# 0.0052f
C268 TEXT$24_0/m3_7680_0# TEXT$8_0/m4_9600_0# 0
C269 TEXT$4_0/m3_8400_0# TEXT$4_0/m3_9600_0# 0.30861f
C270 TEXT$21_0/m4_15120_0# TEXT$7_0/m2_10560_0# 0
C271 TEXT$21_0/m4_4320_0# TEXT$20_0/m3_4320_0# 0.40732f
C272 TEXT$22_0/m2_16560_0# TEXT$21_0/m4_16560_0# 0.0038f
C273 TEXT$24_0/m3_3840_0# TEXT$24_0/m3_4800_960# 0.15024f
C274 TEXT$9_0/m1_10560_0# TEXT$8_0/m4_9600_0# -0
C275 TEXT$7_0/m2_9600_0# TEXT$20_0/m3_14400_0# 0
C276 TEXT$4_0/m3_8400_0# TEXT$6_0/m4_8400_0# 1.13298f
C277 TEXT$22_0/m2_15840_0# TEXT$20_0/m3_15840_0# 0.40709f
C278 TEXT$22_0/m2_15120_0# TEXT$8_0/m4_10560_0# 0
C279 TEXT$22_0/m2_10800_0# TEXT$9_0/m1_6720_0# 0
C280 TEXT$22_0/m2_12960_0# TEXT$3_0/m2_10800_0# 0.00873f
C281 TEXT$21_0/m4_10800_0# TEXT$24_0/m3_6720_0# 0
C282 TEXT$4_0/m3_9600_0# TEXT$3_0/m2_8400_0# 0
C283 TEXT$22_0/m2_4320_0# TEXT$1_0/m1_2400_0# 0
C284 TEXT$3_0/m2_8400_0# TEXT$6_0/m4_8400_0# 0.00893f
C285 TEXT$22_0/m2_15120_0# TEXT$23_0/m1_15120_0# 0.36457f
C286 TEXT$24_0/m3_5760_0# TEXT$9_0/m1_5760_0# 0.01213f
C287 TEXT$7_0/m2_2160_0# VDD 0.0166f
C288 TEXT$21_0/m4_7200_0# TEXT$7_0/m2_2880_0# 0
C289 TEXT$3_0/m2_0_0# TEXT$20_0/m3_2880_720# 0
C290 TEXT$22_0/m2_7200_0# TEXT$23_0/m1_7200_0# 0.36389f
C291 TEXT$1_0/m1_9600_0# TEXT$1_0/m1_10800_0# 0.13176f
C292 TEXT$21_0/m4_13680_0# TEXT$21_0/m4_14400_0# 0.27086f
C293 TEXT$21_0/m4_12960_0# TEXT$20_0/m3_13680_0# 0
C294 TEXT$21_0/m4_10080_0# TEXT$6_0/m4_7200_0# 0.02119f
C295 TEXT$21_0/m4_13680_0# TEXT$20_0/m3_12960_0# 0
C296 TEXT$1_0/m1_6000_0# TEXT$6_0/m4_6000_0# 0.00492f
C297 TEXT$8_0/m4_6720_0# TEXT$20_0/m3_11700_0# 0
C298 TEXT$20_0/m3_11700_0# TEXT$20_0/m3_12960_0# 0.02412f
C299 TEXT$20_0/m3_2880_720# TEXT$20_0/m3_3780_0# 0.09503f
C300 TEXT$6_0/m4_1200_0# TEXT$6_0/m4_2400_0# 0.29078f
C301 TEXT$21_0/m4_0_0# TEXT$20_0/m3_0_0# 0.44276f
C302 TEXT$23_0/m1_14400_0# TEXT$8_0/m4_9600_0# -0
C303 TEXT$22_0/m2_11700_0# TEXT$7_0/m2_7680_0# 0.00282f
C304 TEXT$4_0/m3_2400_0# TEXT$20_0/m3_4320_0# 0.00835f
C305 TEXT$1_0/m1_1200_0# TEXT$3_0/m2_1200_0# 1.11971f
C306 TEXT$8_0/m4_5760_0# VDD 0.00865f
C307 TEXT$21_0/m4_6480_0# TEXT$8_0/m4_2160_0# 0.01474f
C308 TEXT$22_0/m2_10800_0# TEXT$23_0/m1_11700_0# 0
C309 TEXT$24_0/m3_4800_960# TEXT$9_0/m1_3840_0# 0
C310 TEXT$24_0/m3_3840_0# TEXT$9_0/m1_4800_960# 0
C311 TEXT$23_0/m1_7920_720# TEXT$1_0/m1_6000_0# 0.00818f
C312 TEXT$21_0/m4_6480_0# TEXT$22_0/m2_6480_0# 0.004f
C313 TEXT$21_0/m4_11700_0# TEXT$23_0/m1_12960_0# -0
C314 TEXT$1_0/m1_1200_0# TEXT$20_0/m3_4320_0# 0
C315 TEXT$1_0/m1_8400_0# TEXT$23_0/m1_11700_0# 0
C316 TEXT$21_0/m4_12960_0# TEXT$23_0/m1_11700_0# 0
C317 TEXT$23_0/m1_6480_0# TEXT$22_0/m2_5760_0# 0.00148f
C318 TEXT$23_0/m1_10800_0# TEXT$20_0/m3_11700_0# 0
C319 sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# PD 0.00461f
C320 TEXT$22_0/m2_0_0# TEXT$20_0/m3_0_0# 0.44472f
C321 VDD TEXT$7_0/m2_6720_0# 0.0304f
C322 TEXT$21_0/m4_7200_0# TEXT$23_0/m1_6480_0# 0
C323 TEXT$6_0/m4_6000_0# TEXT$20_0/m3_8640_0# 0
C324 TEXT$24_0/m3_0_0# TEXT$23_0/m1_4320_0# 0
C325 TEXT$22_0/m2_5760_0# TEXT$7_0/m2_960_0# 0.00449f
C326 TEXT$22_0/m2_4320_0# TEXT$3_0/m2_2400_0# 0.00513f
C327 TEXT$21_0/m4_6480_0# TEXT$7_0/m2_2160_0# 0
C328 TEXT$22_0/m2_11700_0# TEXT$21_0/m4_10800_0# 0
C329 TEXT$21_0/m4_17280_0# TEXT$23_0/m1_18000_0# -0
C330 TEXT$4_0/m3_10800_0# TEXT$1_0/m1_9600_0# 0.00129f
C331 TEXT$23_0/m1_9360_0# TEXT$22_0/m2_9360_0# 0.41722f
C332 TEXT$21_0/m4_12960_0# TEXT$6_0/m4_10800_0# 0.01349f
C333 TEXT$4_0/m3_6000_0# TEXT$6_0/m4_6000_0# 1.12204f
C334 TEXT$1_0/m1_9600_0# TEXT$6_0/m4_9600_0# 0.00495f
C335 TEXT$8_0/m4_9600_0# VDD 0.01299f
C336 TEXT$6_0/m4_9600_0# TEXT$20_0/m3_11700_0# 0
C337 TEXT$8_0/m4_0_0# TEXT$7_0/m2_960_0# 0
C338 TEXT$22_0/m2_5760_0# TEXT$20_0/m3_4320_0# 0
C339 TEXT$22_0/m2_4320_0# TEXT$20_0/m3_5760_0# 0
C340 TEXT$21_0/m4_4320_0# TEXT$24_0/m3_0_0# 0
C341 TEXT$21_0/m4_5760_0# TEXT$22_0/m2_6480_0# 0
C342 BCM_OUT VDD 0.12526f
C343 TEXT$21_0/m4_6480_0# TEXT$20_0/m3_5760_0# 0.00142f
C344 TEXT$3_0/m2_6000_0# TEXT$6_0/m4_6000_0# 0.0097f
C345 TEXT$4_0/m3_8400_0# TEXT$23_0/m1_11700_0# 0
C346 TEXT$9_0/m1_3840_0# TEXT$9_0/m1_4800_960# 0.11093f
C347 TEXT$8_0/m4_0_0# TEXT$20_0/m3_4320_0# 0
C348 TEXT$22_0/m2_16560_0# TEXT$21_0/m4_17280_0# 0
C349 TEXT$24_0/m3_7680_0# TEXT$7_0/m2_9600_0# 0
C350 TEXT$24_0/m3_9600_0# TEXT$7_0/m2_7680_0# 0
C351 TEXT$23_0/m1_17280_0# TEXT$20_0/m3_17280_0# 0.00325f
C352 TEXT$6_0/m4_6000_0# TEXT$20_0/m3_7920_720# 0
C353 m3_419992_265695# a_498947_268180# 1.74671f
C354 TEXT$9_0/m1_9600_0# TEXT$7_0/m2_10560_0# 0
C355 TEXT$9_0/m1_10560_0# TEXT$7_0/m2_9600_0# 0.00466f
C356 TEXT$23_0/m1_7920_720# TEXT$3_0/m2_6000_0# 0
C357 TEXT$9_0/m1_4800_960# TEXT$9_0/m1_5760_0# 0.12596f
C358 TEXT$24_0/m3_7680_0# TEXT$8_0/m4_7680_0# 0.72108f
C359 TEXT$23_0/m1_15120_0# TEXT$3_0/m2_12000_0# 0
C360 TEXT$21_0/m4_8640_0# TEXT$7_0/m2_3840_0# 0
C361 TEXT$3_0/m2_1200_0# TEXT$20_0/m3_4320_0# 0
C362 TEXT$3_0/m2_8400_0# TEXT$23_0/m1_11700_0# 0
C363 TEXT$23_0/m1_10080_0# TEXT$22_0/m2_9360_0# 0
C364 TEXT$23_0/m1_7920_720# TEXT$20_0/m3_7920_720# 0.00212f
C365 VDD PD 0.05396f
C366 TEXT$24_0/m3_10560_0# TEXT$8_0/m4_9600_0# 0.00399f
C367 TEXT$9_0/m1_5760_0# TEXT$9_0/m1_6720_0# 0.21606f
C368 TEXT$4_0/m3_9600_0# TEXT$4_0/m3_10800_0# 0.16583f
C369 CCM_OUT VDD 0.12526f
C370 TEXT$21_0/m4_5760_0# TEXT$20_0/m3_5760_0# 0.40749f
C371 TEXT$21_0/m4_10800_0# TEXT$23_0/m1_10080_0# 0
C372 TEXT$24_0/m3_960_0# VDD 0.00595f
C373 TEXT$7_0/m2_10560_0# TEXT$20_0/m3_15120_0# 0
C374 TEXT$4_0/m3_9600_0# TEXT$6_0/m4_9600_0# 1.01255f
C375 TEXT$22_0/m2_10800_0# TEXT$24_0/m3_6720_0# 0
C376 TEXT$22_0/m2_16560_0# TEXT$20_0/m3_16560_0# 0.40324f
C377 TEXT$6_0/m4_8400_0# TEXT$6_0/m4_9600_0# 0.31031f
C378 TEXT$23_0/m1_4320_0# TEXT$9_0/m1_0_0# 0.01121f
C379 TEXT$21_0/m4_18000_0# TEXT$20_0/m3_17280_0# 0
C380 TEXT$21_0/m4_11700_0# TEXT$24_0/m3_7680_0# 0
C381 TEXT$9_0/m1_6720_0# TEXT$8_0/m4_6720_0# 0.00178f
C382 TEXT$22_0/m2_5760_0# TEXT$1_0/m1_3600_0# 0
C383 TEXT$9_0/m1_7680_0# TEXT$20_0/m3_11700_0# 0
C384 TEXT$22_0/m2_7200_0# TEXT$7_0/m2_2880_0# 0.02191f
C385 TEXT$23_0/m1_14400_0# TEXT$7_0/m2_9600_0# 0
C386 TEXT$4_0/m3_2400_0# TEXT$4_0/m3_3600_0# 0.23558f
C387 TEXT$22_0/m2_15840_0# TEXT$23_0/m1_15840_0# 0.40272f
C388 TEXT$21_0/m4_7920_720# TEXT$21_0/m4_8640_0# 0.10641f
C389 TEXT$21_0/m4_4320_0# TEXT$9_0/m1_0_0# -0.00116f
C390 TEXT$23_0/m1_6480_0# TEXT$1_0/m1_3600_0# 0.00996f
C391 TEXT$22_0/m2_10080_0# TEXT$6_0/m4_7200_0# 0
C392 TEXT$23_0/m1_8640_0# TEXT$8_0/m4_4800_960# -0
C393 TEXT$21_0/m4_14400_0# TEXT$1_0/m1_12000_0# -0
C394 TEXT$1_0/m1_10800_0# TEXT$1_0/m1_12000_0# 0.13202f
C395 TEXT$21_0/m4_14400_0# TEXT$21_0/m4_15120_0# 0.25667f
C396 TEXT$21_0/m4_14400_0# TEXT$20_0/m3_13680_0# 0
C397 TEXT$1_0/m1_7200_0# TEXT$6_0/m4_7200_0# 0.00392f
C398 TEXT$23_0/m1_10800_0# TEXT$9_0/m1_6720_0# 0.01245f
C399 TEXT$20_0/m3_12960_0# TEXT$20_0/m3_13680_0# 0.20543f
C400 TEXT$22_0/m2_6480_0# TEXT$8_0/m4_2160_0# 0
C401 TEXT$6_0/m4_2400_0# TEXT$6_0/m4_3600_0# 0.24184f
C402 TEXT$1_0/m1_2400_0# TEXT$3_0/m2_2400_0# 1.01384f
C403 TEXT$21_0/m4_7200_0# TEXT$22_0/m2_7200_0# 0.00385f
C404 TEXT$21_0/m4_12960_0# TEXT$23_0/m1_13680_0# -0
C405 TEXT$21_0/m4_13680_0# TEXT$23_0/m1_12960_0# 0
C406 TEXT$23_0/m1_11700_0# TEXT$8_0/m4_6720_0# -0
C407 TEXT$23_0/m1_11700_0# TEXT$20_0/m3_12960_0# 0
C408 TEXT$23_0/m1_12960_0# TEXT$20_0/m3_11700_0# 0
C409 TEXT$4_0/m3_3600_0# TEXT$22_0/m2_5760_0# 0
C410 TEXT$8_0/m4_0_0# TEXT$24_0/m3_0_0# 0.60142f
C411 TEXT$7_0/m2_2160_0# TEXT$8_0/m4_2160_0# 0.00739f
C412 VDD TEXT$7_0/m2_9600_0# 0.0415f
C413 TEXT$22_0/m2_14400_0# TEXT$8_0/m4_9600_0# 0
C414 TEXT$9_0/m1_960_0# VDD 0.03045f
C415 TEXT$6_0/m4_7200_0# TEXT$20_0/m3_9360_0# 0
C416 TEXT$24_0/m3_0_0# TEXT$7_0/m2_960_0# 0
C417 TEXT$24_0/m3_960_0# TEXT$7_0/m2_0_0# 0.00769f
C418 TEXT$22_0/m2_6480_0# TEXT$7_0/m2_2160_0# 0.00963f
C419 TEXT$20_0/m3_7920_720# TEXT$23_0/m1_7200_0# 0
C420 TEXT$22_0/m2_11700_0# TEXT$22_0/m2_10800_0# 0.10044f
C421 TEXT$4_0/m3_3600_0# TEXT$23_0/m1_6480_0# 0
C422 TEXT$8_0/m4_7680_0# VDD 0.0052f
C423 TEXT$22_0/m2_5760_0# TEXT$3_0/m2_3600_0# 0.01126f
C424 VIN_OUT VDD 0.0609f
C425 TEXT$23_0/m1_10800_0# TEXT$23_0/m1_11700_0# 0.10298f
C426 TEXT$22_0/m2_12960_0# TEXT$21_0/m4_11700_0# 0
C427 TEXT$22_0/m2_11700_0# TEXT$1_0/m1_8400_0# 0
C428 TEXT$22_0/m2_11700_0# TEXT$21_0/m4_12960_0# 0
C429 TEXT$4_0/m3_12000_0# TEXT$21_0/m4_14400_0# 0
C430 TEXT$4_0/m3_10800_0# TEXT$1_0/m1_12000_0# 0
C431 TEXT$4_0/m3_12000_0# TEXT$1_0/m1_10800_0# 0.00103f
C432 TEXT$4_0/m3_7200_0# TEXT$6_0/m4_7200_0# 0.65343f
C433 TEXT$1_0/m1_10800_0# TEXT$6_0/m4_10800_0# 0.00425f
C434 TEXT$7_0/m2_4800_960# TEXT$7_0/m2_5760_0# 0.12026f
C435 TEXT$20_0/m3_0_0# TEXT$23_0/m1_0_0# 0.00265f
C436 TEXT$6_0/m4_10800_0# TEXT$20_0/m3_12960_0# 0
C437 TEXT$24_0/m3_0_0# TEXT$20_0/m3_4320_0# 0.01493f
C438 TEXT$22_0/m2_6480_0# TEXT$20_0/m3_5760_0# 0
C439 TEXT$22_0/m2_5760_0# TEXT$20_0/m3_6480_0# 0.00225f
C440 TEXT$21_0/m4_5760_0# TEXT$24_0/m3_960_0# 0
C441 TEXT$23_0/m1_6480_0# TEXT$3_0/m2_3600_0# 0
C442 TEXT$7_0/m2_6720_0# TEXT$20_0/m3_10800_0# 0
C443 TEXT$21_0/m4_7200_0# TEXT$20_0/m3_6480_0# 0
C444 TEXT$21_0/m4_2160_0# TEXT$6_0/m4_0_0# 0.01349f
C445 TEXT$23_0/m1_6480_0# TEXT$20_0/m3_6480_0# 0.00322f
C446 TEXT$24_0/m3_3840_0# TEXT$23_0/m1_7920_720# 0
C447 TEXT$3_0/m2_7200_0# TEXT$6_0/m4_7200_0# 0.00371f
C448 TEXT$24_0/m3_4800_960# TEXT$23_0/m1_8640_0# 0
C449 TEXT$22_0/m2_18000_0# TEXT$21_0/m4_17280_0# 0
C450 TEXT$21_0/m4_8640_0# TEXT$22_0/m2_8640_0# 0.00401f
C451 TEXT$24_0/m3_10560_0# TEXT$7_0/m2_9600_0# 0.00599f
C452 TEXT$24_0/m3_9600_0# TEXT$7_0/m2_10560_0# 0
C453 TEXT$23_0/m1_18000_0# TEXT$20_0/m3_18000_0# 0.00233f
C454 TEXT$4_0/m3_0_0# TEXT$6_0/m4_0_0# 1.13749f
C455 TEXT$22_0/m2_8640_0# TEXT$7_0/m2_3840_0# 0.00481f
C456 TEXT$21_0/m4_9360_0# TEXT$7_0/m2_4800_960# 0
C457 TEXT$8_0/m4_3840_0# TEXT$7_0/m2_2880_0# 0
C458 TEXT$24_0/m3_6720_0# TEXT$9_0/m1_5760_0# 0
C459 TEXT$23_0/m1_10080_0# TEXT$22_0/m2_10800_0# 0
C460 TEXT$21_0/m4_10080_0# TEXT$20_0/m3_10800_0# 0
C461 TEXT$22_0/m2_11700_0# TEXT$4_0/m3_8400_0# 0
C462 TEXT$9_0/m1_6720_0# TEXT$9_0/m1_7680_0# 0.30249f
C463 TEXT$4_0/m3_10800_0# TEXT$4_0/m3_12000_0# 0.14777f
C464 TEXT$8_0/m4_0_0# TEXT$9_0/m1_0_0# 0.00223f
C465 TEXT$22_0/m2_17280_0# TEXT$20_0/m3_17280_0# 0.41033f
C466 TEXT$4_0/m3_10800_0# TEXT$6_0/m4_10800_0# 1.15953f
C467 TEXT$6_0/m4_9600_0# TEXT$6_0/m4_10800_0# 0.17351f
C468 TEXT$8_0/m4_10560_0# TEXT$7_0/m2_10560_0# 0.01523f
C469 TEXT$8_0/m4_2880_0# TEXT$23_0/m1_7200_0# -0.00109f
C470 TEXT$9_0/m1_0_0# TEXT$7_0/m2_960_0# 0
C471 TEXT$9_0/m1_960_0# TEXT$7_0/m2_0_0# 0.00386f
C472 TEXT$22_0/m2_15120_0# TEXT$3_0/m2_12000_0# 0.00625f
C473 TEXT$24_0/m3_6720_0# TEXT$8_0/m4_6720_0# 0.71314f
C474 TEXT$22_0/m2_11700_0# TEXT$3_0/m2_8400_0# 0
C475 TEXT$24_0/m3_7680_0# TEXT$20_0/m3_11700_0# 0.00469f
C476 TEXT$21_0/m4_8640_0# TEXT$22_0/m2_7920_720# 0
C477 TEXT$21_0/m4_14400_0# TEXT$9_0/m1_9600_0# -0.00251f
C478 TEXT$24_0/m3_2880_0# VDD 0.00519f
C479 TEXT$22_0/m2_7920_720# TEXT$7_0/m2_3840_0# 0.00677f
C480 TEXT$23_0/m1_7920_720# TEXT$9_0/m1_3840_0# 0.00617f
C481 TEXT$24_0/m3_2160_0# TEXT$7_0/m2_2880_0# 0
C482 TEXT$23_0/m1_15120_0# TEXT$7_0/m2_10560_0# 0
C483 TEXT$21_0/m4_7920_720# TEXT$1_0/m1_4800_0# 0
C484 TEXT$22_0/m2_16560_0# TEXT$23_0/m1_16560_0# 0.40019f
C485 TEXT$9_0/m1_0_0# TEXT$20_0/m3_4320_0# 0
C486 TEXT$9_0/m1_4800_960# TEXT$23_0/m1_8640_0# 0.00996f
C487 TEXT$21_0/m4_5760_0# TEXT$9_0/m1_960_0# 0
C488 TEXT$21_0/m4_18000_0# TEXT$23_0/m1_17280_0# 0
C489 TEXT$21_0/m4_0_0# TEXT$21_0/m4_720_0# 0.23216f
C490 TEXT$23_0/m1_10080_0# TEXT$20_0/m3_10080_0# 0.00332f
C491 TEXT$4_0/m3_3600_0# TEXT$1_0/m1_3600_0# 0.01216f
C492 TEXT$24_0/m3_6720_0# TEXT$23_0/m1_10800_0# 0
C493 TEXT$21_0/m4_15120_0# TEXT$21_0/m4_15840_0# 0.21282f
C494 TEXT$21_0/m4_15120_0# TEXT$20_0/m3_14400_0# 0.00146f
C495 TEXT$21_0/m4_14400_0# TEXT$20_0/m3_15120_0# 0
C496 TEXT$23_0/m1_11700_0# TEXT$9_0/m1_7680_0# 0.00279f
C497 TEXT$20_0/m3_13680_0# TEXT$20_0/m3_14400_0# 0.26985f
C498 TEXT$6_0/m4_3600_0# TEXT$6_0/m4_4800_0# 0.33857f
C499 TEXT$24_0/m3_960_0# TEXT$8_0/m4_2160_0# 0
C500 TEXT$24_0/m3_2160_0# TEXT$22_0/m2_5760_0# 0
C501 TEXT$22_0/m2_14400_0# TEXT$7_0/m2_9600_0# 0.00658f
C502 TEXT$1_0/m1_3600_0# TEXT$3_0/m2_3600_0# 1.09919f
C503 TEXT$21_0/m4_720_0# TEXT$22_0/m2_0_0# 0
C504 TEXT$21_0/m4_7920_720# TEXT$22_0/m2_7920_720# 0.00246f
C505 TEXT$1_0/m1_3600_0# TEXT$20_0/m3_6480_0# 0
C506 TEXT$21_0/m4_14400_0# TEXT$23_0/m1_13680_0# 0
C507 TEXT$23_0/m1_13680_0# TEXT$20_0/m3_12960_0# 0
C508 TEXT$22_0/m2_2880_720# TEXT$6_0/m4_0_0# 0
C509 TEXT$24_0/m3_2160_0# TEXT$23_0/m1_6480_0# 0
C510 TEXT$21_0/m4_3780_0# TEXT$6_0/m4_1200_0# 0.01128f
C511 TEXT$21_0/m4_10080_0# TEXT$8_0/m4_5760_0# 0.02513f
C512 TEXT$9_0/m1_2880_0# VDD 0.02823f
C513 TEXT$4_0/m3_4800_0# TEXT$21_0/m4_7920_720# 0
C514 TEXT$24_0/m3_960_0# TEXT$7_0/m2_2160_0# 0
C515 TEXT$24_0/m3_2160_0# TEXT$7_0/m2_960_0# 0.00227f
C516 TEXT$24_0/m3_2880_0# TEXT$21_0/m4_6480_0# 0
C517 TEXT$8_0/m4_4800_960# VDD 0.0026f
C518 TEXT$23_0/m1_11700_0# TEXT$23_0/m1_12960_0# 0.0152f
C519 TEXT$22_0/m2_0_0# TEXT$22_0/m2_720_0# 0.19794f
C520 TEXT$22_0/m2_11700_0# TEXT$8_0/m4_6720_0# 0
C521 TEXT$22_0/m2_13680_0# TEXT$21_0/m4_12960_0# 0
C522 TEXT$23_0/m1_2160_0# TEXT$6_0/m4_0_0# 0
C523 TEXT$22_0/m2_12960_0# TEXT$21_0/m4_13680_0# 0
C524 TEXT$22_0/m2_11700_0# TEXT$20_0/m3_12960_0# 0
C525 TEXT$22_0/m2_12960_0# TEXT$20_0/m3_11700_0# 0
C526 TEXT$4_0/m3_12000_0# TEXT$20_0/m3_14400_0# 0.03063f
C527 TEXT$21_0/m4_15120_0# TEXT$6_0/m4_12000_0# 0.01f
C528 TEXT$1_0/m1_12000_0# TEXT$6_0/m4_12000_0# 0.00238f
C529 m4_400150_261569# M_0/a_404041_244568# 0.14584f
C530 m3_419992_265695# m4_400150_261569# 0.10503f
C531 TEXT$21_0/m4_7920_720# TEXT$3_0/m2_4800_0# 0
C532 TEXT$6_0/m4_7200_0# TEXT$6_0/m4_8400_0# 0.13128f
C533 TEXT$9_0/m1_2160_0# TEXT$7_0/m2_2880_0# 0
C534 TEXT$24_0/m3_960_0# TEXT$20_0/m3_5760_0# 0.0059f
C535 TEXT$22_0/m2_6480_0# TEXT$20_0/m3_7200_0# 0.00184f
C536 TEXT$4_0/m3_3600_0# TEXT$3_0/m2_3600_0# 1.09551f
C537 TEXT$21_0/m4_7920_720# TEXT$20_0/m3_7200_0# 0
C538 TEXT$21_0/m4_7200_0# TEXT$20_0/m3_7920_720# 0
C539 TEXT$6_0/m4_0_0# TEXT$20_0/m3_2160_0# 0
C540 TEXT$22_0/m2_11700_0# TEXT$23_0/m1_10800_0# 0
C541 TEXT$4_0/m3_3600_0# TEXT$20_0/m3_6480_0# 0.01525f
C542 TEXT$21_0/m4_9360_0# TEXT$22_0/m2_9360_0# 0.00452f
C543 TEXT$23_0/m1_12960_0# TEXT$6_0/m4_10800_0# 0
C544 TEXT$4_0/m3_1200_0# TEXT$6_0/m4_1200_0# 1.12172f
C545 TEXT$9_0/m1_960_0# TEXT$8_0/m4_2160_0# 0
C546 TEXT$24_0/m3_5760_0# VDD 0.00595f
C547 TEXT$22_0/m2_9360_0# TEXT$7_0/m2_4800_960# 0.01074f
C548 TEXT$23_0/m1_10080_0# TEXT$9_0/m1_5760_0# 0.01607f
C549 TEXT$24_0/m3_0_0# TEXT$9_0/m1_0_0# 0.01017f
C550 TEXT$1_0/m1_1200_0# TEXT$6_0/m4_0_0# 0
C551 TEXT$3_0/m2_3600_0# TEXT$20_0/m3_6480_0# 0
C552 TEXT$22_0/m2_10080_0# TEXT$20_0/m3_10800_0# 0.00285f
C553 TEXT$24_0/m3_7680_0# TEXT$9_0/m1_6720_0# 0
C554 a_498947_268180# a_499016_248165# 0.09669f
C555 TEXT$23_0/m1_6480_0# TEXT$9_0/m1_2160_0# 0.00868f
C556 TEXT$9_0/m1_7680_0# TEXT$9_0/m1_9600_0# 0.02044f
C557 TEXT$8_0/m4_2880_0# TEXT$7_0/m2_2880_0# 0.01326f
C558 TEXT$21_0/m4_11700_0# TEXT$20_0/m3_10800_0# 0
C559 TEXT$22_0/m2_11700_0# TEXT$6_0/m4_9600_0# 0
C560 TEXT$22_0/m2_18000_0# TEXT$20_0/m3_18000_0# 0.34869f
C561 TEXT$4_0/m3_12000_0# TEXT$6_0/m4_12000_0# 1.11712f
C562 TEXT$6_0/m4_10800_0# TEXT$6_0/m4_12000_0# 0.14856f
C563 TEXT$8_0/m4_960_0# VDD 0.00865f
C564 TEXT$22_0/m2_7920_720# TEXT$22_0/m2_8640_0# 0.07523f
C565 TEXT$9_0/m1_960_0# TEXT$7_0/m2_2160_0# 0
C566 TEXT$9_0/m1_2160_0# TEXT$7_0/m2_960_0# 0.00132f
C567 TEXT$21_0/m4_14400_0# TEXT$24_0/m3_9600_0# 0.00155f
C568 TEXT$21_0/m4_15120_0# TEXT$9_0/m1_10560_0# 0
C569 TEXT$22_0/m2_7920_720# TEXT$1_0/m1_4800_0# 0
C570 TEXT$21_0/m4_9360_0# TEXT$20_0/m3_8640_0# 0
C571 TEXT$24_0/m3_4800_960# VDD 0.00195f
C572 TEXT$9_0/m1_9600_0# TEXT$20_0/m3_14400_0# 0
C573 TEXT$22_0/m2_4320_0# TEXT$6_0/m4_1200_0# 0
C574 PU sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# 0.00439f
C575 TEXT$20_0/m3_8640_0# TEXT$7_0/m2_4800_960# 0
C576 TEXT$22_0/m2_17280_0# TEXT$23_0/m1_17280_0# 0.4026f
C577 TEXT$23_0/m1_10080_0# TEXT$23_0/m1_10800_0# 0.27388f
C578 TEXT$9_0/m1_960_0# TEXT$20_0/m3_5760_0# 0
C579 M_0/a_401151_244568# a_498947_268180# 0.01586f
C580 TEXT$21_0/m4_720_0# TEXT$21_0/m4_1440_0# 0.27086f
C581 TEXT$21_0/m4_7200_0# TEXT$8_0/m4_2880_0# 0.03173f
C582 TEXT$4_0/m3_4800_0# TEXT$1_0/m1_4800_0# 0.01052f
C583 TEXT$24_0/m3_7680_0# TEXT$23_0/m1_11700_0# 0
C584 TEXT$21_0/m4_15840_0# TEXT$21_0/m4_16560_0# 0.26312f
C585 TEXT$21_0/m4_15840_0# TEXT$20_0/m3_15120_0# 0
C586 TEXT$24_0/m3_3840_0# TEXT$7_0/m2_2880_0# 0.00485f
C587 TEXT$20_0/m3_14400_0# TEXT$20_0/m3_15120_0# 0.25479f
C588 TEXT$6_0/m4_4800_0# TEXT$6_0/m4_6000_0# 0.26602f
C589 TEXT$21_0/m4_14400_0# TEXT$8_0/m4_10560_0# 0.01115f
C590 TEXT$23_0/m1_4320_0# TEXT$6_0/m4_2400_0# -0
C591 TEXT$23_0/m1_5760_0# TEXT$22_0/m2_4320_0# 0
C592 TEXT$1_0/m1_8400_0# TEXT$3_0/m2_9600_0# 0.00634f
C593 TEXT$22_0/m2_15120_0# TEXT$7_0/m2_10560_0# 0.01841f
C594 TEXT$1_0/m1_4800_0# TEXT$3_0/m2_4800_0# 1.10268f
C595 TEXT$3_0/m2_1200_0# TEXT$6_0/m4_0_0# 0.00123f
C596 TEXT$21_0/m4_6480_0# TEXT$23_0/m1_5760_0# -0
C597 TEXT$22_0/m2_0_0# TEXT$20_0/m3_720_0# 0.00177f
C598 TEXT$22_0/m2_10080_0# TEXT$8_0/m4_5760_0# 0
C599 TEXT$21_0/m4_1440_0# TEXT$22_0/m2_720_0# 0
C600 TEXT$23_0/m1_7920_720# TEXT$6_0/m4_4800_0# 0
C601 TEXT$22_0/m2_17280_0# TEXT$21_0/m4_18000_0# 0
C602 TEXT$8_0/m4_7680_0# TEXT$7_0/m2_6720_0# 0
C603 TEXT$21_0/m4_14400_0# TEXT$23_0/m1_15120_0# -0
C604 TEXT$1_0/m1_12000_0# TEXT$23_0/m1_14400_0# 0.01915f
C605 TEXT$21_0/m4_15120_0# TEXT$23_0/m1_14400_0# 0
C606 TEXT$24_0/m3_2880_0# TEXT$8_0/m4_2160_0# 0.00169f
C607 TEXT$6_0/m4_1200_0# TEXT$20_0/m3_3780_0# 0
C608 TEXT$6_0/m4_6000_0# TEXT$23_0/m1_8640_0# -0
C609 TEXT$22_0/m2_11700_0# TEXT$9_0/m1_7680_0# 0
C610 TEXT$21_0/m4_4320_0# TEXT$6_0/m4_2400_0# 0.00842f
C611 TEXT$24_0/m3_2880_0# TEXT$22_0/m2_6480_0# 0
C612 TEXT$4_0/m3_4800_0# TEXT$22_0/m2_7920_720# 0
C613 TEXT$8_0/m4_9600_0# TEXT$7_0/m2_9600_0# 0.01727f
C614 TEXT$9_0/m1_4800_960# VDD 0.00782f
C615 m4_400150_261569# a_498947_268180# 0.07748f
C616 TEXT$23_0/m1_7920_720# TEXT$23_0/m1_8640_0# 0.07639f
C617 TEXT$8_0/m4_960_0# TEXT$7_0/m2_0_0# 0
C618 TEXT$21_0/m4_720_0# TEXT$23_0/m1_0_0# 0
C619 TEXT$8_0/m4_7680_0# TEXT$8_0/m4_9600_0# 0.03495f
C620 TEXT$22_0/m2_7920_720# TEXT$3_0/m2_4800_0# 0.00794f
C621 VDD VBIAS 19.64782f
C622 TEXT$23_0/m1_12960_0# TEXT$23_0/m1_13680_0# 0.22968f
C623 TEXT$21_0/m4_11700_0# TEXT$7_0/m2_6720_0# 0
C624 TEXT$9_0/m1_6720_0# VDD 0.03281f
C625 TEXT$22_0/m2_13680_0# TEXT$21_0/m4_14400_0# 0
C626 TEXT$22_0/m2_13680_0# TEXT$20_0/m3_12960_0# 0
C627 TEXT$22_0/m2_12960_0# TEXT$20_0/m3_13680_0# 0.00261f
C628 TEXT$22_0/m2_7920_720# TEXT$20_0/m3_7200_0# 0
C629 TEXT$22_0/m2_7200_0# TEXT$20_0/m3_7920_720# 0.00101f
C630 TEXT$6_0/m4_12000_0# TEXT$20_0/m3_15120_0# 0
C631 TEXT$24_0/m3_2880_0# TEXT$7_0/m2_2160_0# 0.00228f
C632 TEXT$9_0/m1_2880_0# TEXT$7_0/m2_3840_0# 0.00137f
C633 TEXT$9_0/m1_3840_0# TEXT$7_0/m2_2880_0# 0.00209f
C634 TEXT$24_0/m3_2160_0# TEXT$20_0/m3_6480_0# 0.01353f
C635 TEXT$23_0/m1_720_0# TEXT$22_0/m2_0_0# 0.00159f
C636 TEXT$21_0/m4_5760_0# TEXT$23_0/m1_5760_0# -0
C637 TEXT$21_0/m4_8640_0# TEXT$8_0/m4_4800_960# 0.01644f
C638 TEXT$22_0/m2_3780_0# TEXT$23_0/m1_3780_0# 0.19314f
C639 TEXT$4_0/m3_8400_0# TEXT$3_0/m2_9600_0# 0
C640 TEXT$8_0/m4_4800_960# TEXT$7_0/m2_3840_0# 0
C641 TEXT$8_0/m4_960_0# TEXT$21_0/m4_5760_0# 0.00683f
C642 TEXT$4_0/m3_4800_0# TEXT$3_0/m2_4800_0# 1.09377f
C643 TEXT$4_0/m3_4800_0# TEXT$20_0/m3_7200_0# 0.02525f
C644 TEXT$22_0/m2_11700_0# TEXT$23_0/m1_12960_0# 0
C645 TEXT$22_0/m2_12960_0# TEXT$23_0/m1_11700_0# 0
C646 TEXT$21_0/m4_10080_0# TEXT$22_0/m2_10080_0# 0.00591f
C647 TEXT$4_0/m3_2400_0# TEXT$6_0/m4_2400_0# 1.01621f
C648 TEXT$3_0/m2_8400_0# TEXT$3_0/m2_9600_0# 0.24273f
C649 TEXT$9_0/m1_2880_0# TEXT$8_0/m4_2160_0# 0
C650 TEXT$20_0/m3_10080_0# TEXT$7_0/m2_5760_0# 0.00106f
C651 TEXT$21_0/m4_10080_0# TEXT$1_0/m1_7200_0# 0
C652 TEXT$23_0/m1_4320_0# TEXT$23_0/m1_3780_0# 0.10298f
C653 TEXT$23_0/m1_9360_0# TEXT$23_0/m1_8640_0# 0.29377f
C654 TEXT$24_0/m3_960_0# TEXT$9_0/m1_960_0# 0.01213f
C655 TEXT$1_0/m1_1200_0# TEXT$6_0/m4_2400_0# -0.01711f
C656 TEXT$1_0/m1_2400_0# TEXT$6_0/m4_1200_0# 0
C657 TEXT$21_0/m4_1440_0# TEXT$22_0/m2_1440_0# 0.0049f
C658 TEXT$3_0/m2_4800_0# TEXT$20_0/m3_7200_0# 0
C659 TEXT$24_0/m3_6720_0# TEXT$24_0/m3_7680_0# 0.30445f
C660 TEXT$24_0/m3_9600_0# TEXT$9_0/m1_7680_0# 0
C661 TEXT$24_0/m3_7680_0# TEXT$9_0/m1_9600_0# 0
C662 TEXT$9_0/m1_9600_0# TEXT$9_0/m1_10560_0# 0.16595f
C663 TEXT$22_0/m2_3780_0# TEXT$23_0/m1_2880_720# 0
C664 TEXT$22_0/m2_2880_720# TEXT$23_0/m1_3780_0# 0
C665 TEXT$22_0/m2_12960_0# TEXT$6_0/m4_10800_0# 0
C666 TEXT$20_0/m3_10800_0# TEXT$20_0/m3_11700_0# 0.13459f
C667 TEXT$6_0/m4_4800_0# TEXT$23_0/m1_7200_0# 0
C668 TEXT$21_0/m4_4320_0# TEXT$23_0/m1_3780_0# 0
C669 TEXT$9_0/m1_2880_0# TEXT$7_0/m2_2160_0# 0.00129f
C670 TEXT$22_0/m2_8640_0# TEXT$20_0/m3_9360_0# 0.00184f
C671 TEXT$21_0/m4_15120_0# TEXT$24_0/m3_10560_0# 0
C672 TEXT$24_0/m3_9600_0# TEXT$20_0/m3_14400_0# 0.01497f
C673 TEXT$21_0/m4_10080_0# TEXT$20_0/m3_9360_0# 0.00136f
C674 TEXT$8_0/m4_3840_0# TEXT$20_0/m3_8640_0# 0
C675 TEXT$9_0/m1_10560_0# TEXT$20_0/m3_15120_0# 0
C676 TEXT$22_0/m2_18000_0# TEXT$23_0/m1_18000_0# 0.34645f
C677 TEXT$22_0/m2_7200_0# TEXT$8_0/m4_2880_0# 0
C678 TEXT$9_0/m1_2160_0# TEXT$20_0/m3_6480_0# 0
C679 TEXT$21_0/m4_6480_0# TEXT$6_0/m4_3600_0# 0.01714f
C680 TEXT$21_0/m4_1440_0# TEXT$20_0/m3_720_0# 0
C681 TEXT$4_0/m3_7200_0# TEXT$21_0/m4_10080_0# 0
C682 TEXT$4_0/m3_6000_0# TEXT$1_0/m1_6000_0# 0.01243f
C683 TEXT$21_0/m4_1440_0# TEXT$21_0/m4_2160_0# 0.14833f
C684 TEXT$24_0/m3_4800_960# TEXT$21_0/m4_8640_0# 0
C685 TEXT$21_0/m4_16560_0# TEXT$20_0/m3_15840_0# 0
C686 TEXT$24_0/m3_4800_960# TEXT$7_0/m2_3840_0# 0.00319f
C687 TEXT$24_0/m3_3840_0# TEXT$7_0/m2_4800_960# 0
C688 TEXT$23_0/m1_14400_0# TEXT$9_0/m1_9600_0# 0.00972f
C689 TEXT$22_0/m2_2880_720# TEXT$23_0/m1_2880_720# 0.23534f
C690 TEXT$20_0/m3_15120_0# TEXT$20_0/m3_15840_0# 0.22404f
C691 TEXT$6_0/m4_6000_0# TEXT$6_0/m4_7200_0# 0.32706f
C692 TEXT$8_0/m4_4800_960# TEXT$8_0/m4_5760_0# 0.16804f
C693 TEXT$8_0/m4_10560_0# TEXT$20_0/m3_14400_0# 0.00211f
C694 TEXT$23_0/m1_5760_0# TEXT$22_0/m2_6480_0# 0
C695 TEXT$1_0/m1_10800_0# TEXT$3_0/m2_9600_0# 0
C696 TEXT$1_0/m1_9600_0# TEXT$3_0/m2_10800_0# 0.00282f
C697 TEXT$8_0/m4_960_0# TEXT$8_0/m4_2160_0# 0.15081f
C698 TEXT$21_0/m4_10080_0# TEXT$3_0/m2_7200_0# 0
C699 TEXT$1_0/m1_6000_0# TEXT$3_0/m2_6000_0# 1.11971f
C700 TEXT$6_0/m4_8400_0# TEXT$20_0/m3_10800_0# 0
C701 TEXT$3_0/m2_2400_0# TEXT$6_0/m4_1200_0# 0.0019f
C702 TEXT$22_0/m2_720_0# TEXT$20_0/m3_1440_0# 0.0018f
C703 TEXT$21_0/m4_15840_0# TEXT$23_0/m1_15120_0# 0
C704 TEXT$1_0/m1_6000_0# TEXT$20_0/m3_7920_720# 0
C705 TEXT$8_0/m4_3840_0# TEXT$20_0/m3_7920_720# 0
C706 TEXT$22_0/m2_11700_0# TEXT$24_0/m3_7680_0# 0
C707 TEXT$23_0/m1_15120_0# TEXT$20_0/m3_14400_0# 0
C708 TEXT$6_0/m4_2400_0# TEXT$20_0/m3_4320_0# 0
C709 TEXT$21_0/m4_5760_0# TEXT$6_0/m4_3600_0# 0.0166f
C710 TEXT$1_0/m1_1200_0# TEXT$23_0/m1_3780_0# 0.00639f
C711 TEXT$9_0/m1_5760_0# TEXT$7_0/m2_5760_0# 0.65326f
C712 TEXT$23_0/m1_2160_0# TEXT$23_0/m1_2880_720# 0.12753f
C713 TEXT$21_0/m4_1440_0# TEXT$23_0/m1_720_0# 0
C714 TEXT$4_0/m3_6000_0# TEXT$20_0/m3_8640_0# 0.0208f
C715 TEXT$24_0/m3_5760_0# TEXT$8_0/m4_5760_0# 0.66257f
C716 TEXT$22_0/m2_1440_0# TEXT$22_0/m2_2160_0# 0.11417f
C717 TEXT$24_0/m3_6720_0# VDD 0.00864f
C718 TEXT$23_0/m1_13680_0# TEXT$23_0/m1_14400_0# 0.30936f
C719 TEXT$3_0/m2_6000_0# TEXT$20_0/m3_8640_0# 0
C720 TEXT$8_0/m4_6720_0# TEXT$7_0/m2_5760_0# 0
C721 TEXT$9_0/m1_9600_0# VDD 0.03879f
C722 TEXT$22_0/m2_8640_0# TEXT$8_0/m4_4800_960# 0
C723 TEXT$7_0/m2_6720_0# TEXT$20_0/m3_11700_0# 0
C724 TEXT$22_0/m2_14400_0# TEXT$1_0/m1_12000_0# 0
C725 TEXT$22_0/m2_14400_0# TEXT$21_0/m4_15120_0# 0
C726 TEXT$21_0/m4_8640_0# TEXT$9_0/m1_4800_960# 0
C727 TEXT$22_0/m2_13680_0# TEXT$20_0/m3_14400_0# 0.0018f
C728 TEXT$23_0/m1_5760_0# TEXT$20_0/m3_5760_0# 0.00325f
C729 TEXT$9_0/m1_4800_960# TEXT$7_0/m2_3840_0# 0.00247f
C730 TEXT$20_0/m3_7920_720# TEXT$20_0/m3_8640_0# 0.1014f
C731 TEXT$21_0/m4_11700_0# TEXT$8_0/m4_7680_0# 0.00429f
C732 TEXT$8_0/m4_960_0# TEXT$20_0/m3_5760_0# 0
C733 TEXT$23_0/m1_9360_0# TEXT$6_0/m4_7200_0# -0
C734 TEXT$4_0/m3_9600_0# TEXT$3_0/m2_10800_0# 0
C735 TEXT$4_0/m3_10800_0# TEXT$3_0/m2_9600_0# 0
C736 TEXT$4_0/m3_6000_0# TEXT$3_0/m2_6000_0# 1.11291f
C737 TEXT$6_0/m4_9600_0# TEXT$3_0/m2_9600_0# 0.00769f
C738 TEXT$9_0/m1_5760_0# TEXT$7_0/m2_4800_960# 0.00169f
C739 TEXT$21_0/m4_13680_0# TEXT$8_0/m4_9600_0# 0.02016f
C740 TEXT$22_0/m2_13680_0# TEXT$23_0/m1_12960_0# 0
C741 TEXT$21_0/m4_1440_0# TEXT$23_0/m1_1440_0# 0
C742 TEXT$22_0/m2_12960_0# TEXT$23_0/m1_13680_0# 0.00175f
C743 TEXT$4_0/m3_6000_0# TEXT$20_0/m3_7920_720# 0.01319f
C744 TEXT$24_0/m3_2880_0# TEXT$20_0/m3_7200_0# 0.03303f
C745 TEXT$23_0/m1_15120_0# TEXT$6_0/m4_12000_0# 0
C746 TEXT$22_0/m2_10080_0# TEXT$1_0/m1_7200_0# 0
C747 TEXT$21_0/m4_10800_0# TEXT$22_0/m2_10800_0# 0.00342f
C748 TEXT$9_0/m1_6720_0# TEXT$20_0/m3_10800_0# 0
C749 TEXT$23_0/m1_720_0# TEXT$23_0/m1_0_0# 0.26517f
C750 TEXT$21_0/m4_10800_0# TEXT$1_0/m1_8400_0# 0
C751 TEXT$24_0/m3_2160_0# TEXT$9_0/m1_2160_0# 0.00619f
C752 TEXT$22_0/m2_1440_0# TEXT$20_0/m3_1440_0# 0.36906f
C753 TEXT$21_0/m4_2160_0# TEXT$22_0/m2_2160_0# 0.00375f
C754 TEXT$1_0/m1_3600_0# TEXT$6_0/m4_2400_0# 0
C755 TEXT$3_0/m2_6000_0# TEXT$20_0/m3_7920_720# 0
C756 TEXT$24_0/m3_7680_0# TEXT$24_0/m3_9600_0# 0.03244f
C757 TEXT$3_0/m2_1200_0# TEXT$23_0/m1_3780_0# 0
C758 TEXT$24_0/m3_9600_0# TEXT$9_0/m1_10560_0# 0
C759 TEXT$24_0/m3_10560_0# TEXT$9_0/m1_9600_0# 0
C760 TEXT$24_0/m3_5760_0# TEXT$21_0/m4_10080_0# 0
C761 TEXT$8_0/m4_2880_0# TEXT$8_0/m4_3840_0# 0.15093f
C762 TEXT$4_0/m3_0_0# TEXT$22_0/m2_2160_0# 0
C763 TEXT$22_0/m2_11700_0# TEXT$22_0/m2_12960_0# 0.01663f
C764 TEXT$22_0/m2_14400_0# TEXT$4_0/m3_12000_0# 0
C765 TEXT$23_0/m1_10080_0# TEXT$6_0/m4_7200_0# 0
C766 TEXT$22_0/m2_10080_0# TEXT$20_0/m3_9360_0# 0
C767 TEXT$22_0/m2_9360_0# TEXT$20_0/m3_10080_0# 0
C768 TEXT$24_0/m3_10560_0# TEXT$20_0/m3_15120_0# 0.02643f
C769 TEXT$21_0/m4_10800_0# TEXT$20_0/m3_10080_0# 0.00114f
C770 TEXT$22_0/m2_6480_0# TEXT$6_0/m4_3600_0# 0
C771 TEXT$23_0/m1_11700_0# TEXT$20_0/m3_10800_0# 0
C772 TEXT$8_0/m4_10560_0# TEXT$9_0/m1_10560_0# 0.00472f
C773 TEXT$24_0/m3_2160_0# TEXT$8_0/m4_2880_0# 0
C774 TEXT$24_0/m3_4800_960# TEXT$22_0/m2_8640_0# 0
C775 TEXT$4_0/m3_7200_0# TEXT$22_0/m2_10080_0# 0
C776 TEXT$9_0/m1_2880_0# TEXT$20_0/m3_7200_0# 0
C777 TEXT$21_0/m4_7200_0# TEXT$6_0/m4_4800_0# 0.02793f
C778 TEXT$20_0/m3_720_0# TEXT$20_0/m3_1440_0# 0.26985f
C779 TEXT$21_0/m4_1440_0# TEXT$20_0/m3_2160_0# 0
C780 TEXT$21_0/m4_2160_0# TEXT$20_0/m3_1440_0# 0
C781 TEXT$4_0/m3_8400_0# TEXT$21_0/m4_10800_0# 0
C782 TEXT$4_0/m3_7200_0# TEXT$1_0/m1_7200_0# 0.00633f
C783 TEXT$21_0/m4_2160_0# TEXT$21_0/m4_2880_720# 0.15478f
C784 TEXT$24_0/m3_3840_0# TEXT$8_0/m4_3840_0# 0.73416f
C785 TEXT$24_0/m3_9600_0# TEXT$23_0/m1_14400_0# 0
C786 TEXT$4_0/m3_3600_0# TEXT$6_0/m4_2400_0# 0.00637f
C787 TEXT$21_0/m4_16560_0# TEXT$20_0/m3_17280_0# 0
C788 TEXT$23_0/m1_15120_0# TEXT$9_0/m1_10560_0# 0.01663f
C789 TEXT$4_0/m3_0_0# TEXT$21_0/m4_2880_720# 0
C790 TEXT$22_0/m2_10080_0# TEXT$3_0/m2_7200_0# 0.01318f
C791 TEXT$20_0/m3_15840_0# TEXT$20_0/m3_16560_0# 0.26159f
C792 TEXT$21_0/m4_3780_0# TEXT$22_0/m2_3780_0# 0.00207f
C793 TEXT$24_0/m3_960_0# TEXT$23_0/m1_5760_0# 0
C794 TEXT$21_0/m4_14400_0# TEXT$3_0/m2_12000_0# 0
C795 TEXT$1_0/m1_12000_0# TEXT$3_0/m2_10800_0# 0
C796 TEXT$1_0/m1_10800_0# TEXT$3_0/m2_12000_0# 0.00298f
C797 TEXT$4_0/m3_0_0# TEXT$4_0/m3_1200_0# 0.25914f
C798 TEXT$21_0/m4_10800_0# TEXT$3_0/m2_8400_0# 0
C799 TEXT$1_0/m1_7200_0# TEXT$3_0/m2_7200_0# 0.65242f
C800 TEXT$3_0/m2_3600_0# TEXT$6_0/m4_2400_0# 0.00112f
C801 TEXT$8_0/m4_960_0# TEXT$24_0/m3_960_0# 0.66257f
C802 TEXT$21_0/m4_16560_0# TEXT$23_0/m1_15840_0# 0
C803 TEXT$4_0/m3_0_0# TEXT$1_0/m1_0_0# 0.011f
C804 TEXT$6_0/m4_3600_0# TEXT$20_0/m3_5760_0# 0
C805 TEXT$9_0/m1_6720_0# TEXT$7_0/m2_6720_0# 0.70441f
C806 TEXT$22_0/m2_14400_0# TEXT$9_0/m1_9600_0# 0.00133f
C807 TEXT$23_0/m1_1440_0# TEXT$22_0/m2_2160_0# 0
C808 TEXT$8_0/m4_10560_0# TEXT$23_0/m1_14400_0# -0.00209f
C809 TEXT$4_0/m3_7200_0# TEXT$20_0/m3_9360_0# 0.0285f
C810 TEXT$24_0/m3_3840_0# TEXT$20_0/m3_8640_0# 0.01353f
C811 TEXT$22_0/m2_8640_0# TEXT$9_0/m1_4800_960# 0
C812 TEXT$22_0/m2_2160_0# TEXT$22_0/m2_2880_720# 0.11506f
C813 TEXT$24_0/m3_9600_0# VDD 0.00918f
C814 TEXT$23_0/m1_14400_0# TEXT$23_0/m1_15120_0# 0.28224f
C815 TEXT$21_0/m4_2880_720# TEXT$22_0/m2_3780_0# 0
C816 TEXT$22_0/m2_15120_0# TEXT$21_0/m4_15840_0# 0
C817 TEXT$21_0/m4_3780_0# TEXT$22_0/m2_2880_720# 0
C818 TEXT$3_0/m2_7200_0# TEXT$20_0/m3_9360_0# 0
C819 TEXT$22_0/m2_15120_0# TEXT$20_0/m3_14400_0# 0
C820 TEXT$22_0/m2_14400_0# TEXT$20_0/m3_15120_0# 0.00219f
C821 TEXT$21_0/m4_3780_0# TEXT$21_0/m4_4320_0# 0.14096f
C822 TEXT$9_0/m1_3840_0# TEXT$8_0/m4_3840_0# 0.00257f
C823 TEXT$4_0/m3_1200_0# TEXT$22_0/m2_3780_0# 0
C824 TEXT$8_0/m4_7680_0# TEXT$20_0/m3_11700_0# 0
C825 TEXT$4_0/m3_12000_0# TEXT$3_0/m2_10800_0# 0
C826 TEXT$4_0/m3_7200_0# TEXT$3_0/m2_7200_0# 0.65046f
C827 TEXT$6_0/m4_10800_0# TEXT$3_0/m2_10800_0# 0.00864f
C828 TEXT$23_0/m1_2160_0# TEXT$22_0/m2_2160_0# 0.39981f
C829 TEXT$23_0/m1_11700_0# TEXT$7_0/m2_6720_0# 0
C830 TEXT$23_0/m1_1440_0# TEXT$20_0/m3_1440_0# 0.00368f
C831 TEXT$8_0/m4_9600_0# TEXT$20_0/m3_13680_0# 0.00214f
C832 TEXT$22_0/m2_13680_0# TEXT$23_0/m1_14400_0# 0.00168f
C833 TEXT$24_0/m3_3840_0# TEXT$20_0/m3_7920_720# 0.0104f
C834 TEXT$8_0/m4_10560_0# VDD 0.01063f
C835 TEXT$24_0/m3_6720_0# TEXT$20_0/m3_10800_0# 0.02009f
C836 TEXT$22_0/m2_10800_0# TEXT$1_0/m1_8400_0# 0
C837 TEXT$21_0/m4_2160_0# TEXT$3_0/m2_0_0# 0
C838 TEXT$4_0/m3_1200_0# TEXT$23_0/m1_4320_0# 0
C839 TEXT$23_0/m1_5760_0# TEXT$9_0/m1_960_0# 0.00395f
C840 TEXT$21_0/m4_10800_0# TEXT$8_0/m4_6720_0# 0.02077f
C841 TEXT$9_0/m1_3840_0# TEXT$20_0/m3_8640_0# 0
C842 TEXT$24_0/m3_5760_0# TEXT$22_0/m2_10080_0# 0
C843 TEXT$22_0/m2_2160_0# TEXT$20_0/m3_2160_0# 0.40205f
C844 TEXT$21_0/m4_11700_0# TEXT$20_0/m3_11700_0# 0.19343f
C845 TEXT$1_0/m1_4800_0# TEXT$6_0/m4_3600_0# 0
C846 TEXT$21_0/m4_8640_0# TEXT$6_0/m4_6000_0# 0.02105f
C847 TEXT$21_0/m4_2880_720# TEXT$22_0/m2_2880_720# 0.00246f
C848 TEXT$4_0/m3_0_0# TEXT$3_0/m2_0_0# 1.12433f
C849 TEXT$8_0/m4_960_0# TEXT$9_0/m1_960_0# 0.00251f
C850 TEXT$24_0/m3_9600_0# TEXT$24_0/m3_10560_0# 0.17494f
C851 TEXT$8_0/m4_4800_960# TEXT$20_0/m3_9360_0# 0
C852 TEXT$22_0/m2_12960_0# TEXT$22_0/m2_13680_0# 0.17402f
C853 TEXT$22_0/m2_3780_0# TEXT$22_0/m2_4320_0# 0.10044f
C854 TEXT$4_0/m3_1200_0# TEXT$21_0/m4_4320_0# 0
C855 TEXT$22_0/m2_15120_0# TEXT$6_0/m4_12000_0# 0
C856 TEXT$24_0/m3_2880_0# TEXT$9_0/m1_2880_0# 0.01143f
C857 TEXT$21_0/m4_8640_0# TEXT$23_0/m1_7920_720# 0
C858 TEXT$22_0/m2_2880_720# TEXT$1_0/m1_0_0# 0
C859 TEXT$23_0/m1_7920_720# TEXT$7_0/m2_3840_0# 0
C860 TEXT$21_0/m4_10800_0# TEXT$23_0/m1_10800_0# 0
C861 TEXT$21_0/m4_9360_0# TEXT$23_0/m1_8640_0# 0
C862 TEXT$22_0/m2_10800_0# TEXT$20_0/m3_10080_0# 0
C863 TEXT$21_0/m4_3780_0# TEXT$1_0/m1_1200_0# 0
C864 TEXT$23_0/m1_2160_0# TEXT$20_0/m3_1440_0# 0
C865 TEXT$21_0/m4_17280_0# TEXT$20_0/m3_17280_0# 0.40733f
C866 TEXT$23_0/m1_8640_0# TEXT$7_0/m2_4800_960# 0
C867 TEXT$21_0/m4_2880_720# TEXT$23_0/m1_2160_0# 0
C868 TEXT$8_0/m4_10560_0# TEXT$24_0/m3_10560_0# 0.75618f
C869 TEXT$22_0/m2_7200_0# TEXT$6_0/m4_4800_0# 0
C870 TEXT$23_0/m1_4320_0# TEXT$22_0/m2_4320_0# 0.40655f
C871 TEXT$4_0/m3_8400_0# TEXT$22_0/m2_10800_0# 0
C872 TEXT$9_0/m1_3840_0# TEXT$20_0/m3_7920_720# 0
C873 TEXT$24_0/m3_5760_0# TEXT$20_0/m3_9360_0# 0
C874 TEXT$21_0/m4_7920_720# TEXT$6_0/m4_6000_0# 0.01378f
C875 TEXT$20_0/m3_1440_0# TEXT$20_0/m3_2160_0# 0.144f
C876 TEXT$23_0/m1_2160_0# TEXT$1_0/m1_0_0# 0.00794f
C877 TEXT$21_0/m4_2880_720# TEXT$20_0/m3_2160_0# 0
C878 TEXT$21_0/m4_2160_0# TEXT$20_0/m3_2880_720# 0
C879 TEXT$4_0/m3_9600_0# TEXT$21_0/m4_11700_0# 0
C880 TEXT$4_0/m3_8400_0# TEXT$1_0/m1_8400_0# 0.01243f
C881 TEXT$24_0/m3_10560_0# TEXT$23_0/m1_15120_0# 0
C882 TEXT$1_0/m1_7200_0# TEXT$6_0/m4_8400_0# 0
C883 TEXT$21_0/m4_11700_0# TEXT$6_0/m4_8400_0# 0
C884 TEXT$4_0/m3_4800_0# TEXT$6_0/m4_3600_0# 0.01007f
C885 TEXT$4_0/m3_0_0# TEXT$20_0/m3_2880_720# 0.0125f
C886 TEXT$22_0/m2_3780_0# TEXT$20_0/m3_3780_0# 0.1943f
C887 TEXT$22_0/m2_10800_0# TEXT$3_0/m2_8400_0# 0.02223f
C888 TEXT$20_0/m3_16560_0# TEXT$20_0/m3_17280_0# 0.12171f
C889 TEXT$24_0/m3_3840_0# TEXT$8_0/m4_2880_0# 0.00481f
C890 TEXT$24_0/m3_6720_0# TEXT$8_0/m4_5760_0# 0.00499f
C891 TEXT$21_0/m4_4320_0# TEXT$22_0/m2_4320_0# 0.0042f
C892 TEXT$21_0/m4_7920_720# TEXT$23_0/m1_7920_720# 0
C893 PU sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# 0
C894 TEXT$23_0/m1_4320_0# TEXT$7_0/m2_0_0# 0
C895 TEXT$22_0/m2_11700_0# TEXT$20_0/m3_10800_0# 0
C896 TEXT$1_0/m1_0_0# TEXT$20_0/m3_2160_0# 0
C897 TEXT$4_0/m3_1200_0# TEXT$4_0/m3_2400_0# 0.31804f
C898 TEXT$20_0/m3_14400_0# TEXT$3_0/m2_12000_0# 0
C899 TEXT$1_0/m1_8400_0# TEXT$3_0/m2_8400_0# 1.1315f
C900 TEXT$3_0/m2_4800_0# TEXT$6_0/m4_3600_0# 0.00201f
C901 VDD M_0/a_404041_244568# -0.01288f
C902 VDD TEXT$7_0/m2_2880_0# 0.02762f
C903 m3_419992_265695# VDD 1.36032f
C904 TEXT$21_0/m4_16560_0# TEXT$23_0/m1_17280_0# -0
C905 TEXT$4_0/m3_1200_0# TEXT$1_0/m1_1200_0# 0.01243f
C906 TEXT$24_0/m3_6720_0# TEXT$7_0/m2_6720_0# 0.71217f
C907 TEXT$22_0/m2_14400_0# TEXT$24_0/m3_9600_0# 0.00111f
C908 TEXT$9_0/m1_7680_0# TEXT$7_0/m2_7680_0# 0.71495f
C909 TEXT$22_0/m2_15120_0# TEXT$9_0/m1_10560_0# 0
C910 TEXT$23_0/m1_4320_0# TEXT$20_0/m3_3780_0# 0
C911 TEXT$21_0/m4_5760_0# TEXT$23_0/m1_4320_0# 0
C912 TEXT$21_0/m4_4320_0# TEXT$7_0/m2_0_0# 0
C913 TEXT$24_0/m3_4800_960# TEXT$20_0/m3_9360_0# 0.01562f
C914 TEXT$1_0/m1_0_0# TEXT$1_0/m1_1200_0# 0.23454f
C915 TEXT$22_0/m2_2880_720# TEXT$3_0/m2_0_0# 0.00873f
C916 TEXT$21_0/m4_3780_0# TEXT$3_0/m2_1200_0# 0
C917 TEXT$22_0/m2_2880_720# TEXT$20_0/m3_3780_0# 0
C918 TEXT$22_0/m2_3780_0# TEXT$20_0/m3_2880_720# 0
C919 TEXT$23_0/m1_15120_0# TEXT$23_0/m1_15840_0# 0.24307f
C920 TEXT$21_0/m4_14400_0# TEXT$7_0/m2_10560_0# 0
C921 TEXT$21_0/m4_3780_0# TEXT$20_0/m3_4320_0# 0
C922 TEXT$21_0/m4_4320_0# TEXT$20_0/m3_3780_0# 0
C923 TEXT$22_0/m2_15840_0# TEXT$21_0/m4_16560_0# 0
C924 TEXT$7_0/m2_9600_0# TEXT$20_0/m3_13680_0# 0.00166f
C925 TEXT$9_0/m1_9600_0# TEXT$8_0/m4_9600_0# 0.00468f
C926 TEXT$22_0/m2_15120_0# TEXT$20_0/m3_15840_0# 0.00141f
C927 TEXT$21_0/m4_4320_0# TEXT$21_0/m4_5760_0# 0.03386f
C928 TEXT$22_0/m2_14400_0# TEXT$8_0/m4_10560_0# 0
C929 TEXT$4_0/m3_2400_0# TEXT$22_0/m2_4320_0# 0
C930 TEXT$9_0/m1_3840_0# TEXT$8_0/m4_2880_0# 0
C931 TEXT$23_0/m1_2160_0# TEXT$3_0/m2_0_0# 0
C932 VDD M_0/a_403251_244568# -0.01121f
C933 TEXT$4_0/m3_8400_0# TEXT$3_0/m2_8400_0# 1.12534f
C934 TEXT$6_0/m4_12000_0# TEXT$3_0/m2_12000_0# 0.01086f
C935 TEXT$21_0/m4_11700_0# TEXT$9_0/m1_6720_0# -0
C936 TEXT$22_0/m2_4320_0# TEXT$1_0/m1_1200_0# 0
C937 TEXT$8_0/m4_0_0# VDD 0.01058f
C938 TEXT$24_0/m3_5760_0# TEXT$8_0/m4_4800_960# 0.00313f
C939 PU EN 0.21991f
C940 TEXT$22_0/m2_15120_0# TEXT$23_0/m1_14400_0# 0
C941 TEXT$22_0/m2_14400_0# TEXT$23_0/m1_15120_0# 0.00177f
C942 TEXT$7_0/m2_960_0# VDD 0.03306f
C943 TEXT$22_0/m2_10800_0# TEXT$8_0/m4_6720_0# 0
C944 TEXT$3_0/m2_0_0# TEXT$20_0/m3_2160_0# 0
C945 TEXT$22_0/m2_8640_0# TEXT$6_0/m4_6000_0# 0
C946 PU VDD 0.00886f
C947 TEXT$22_0/m2_6480_0# TEXT$23_0/m1_7200_0# 0.00171f
C948 TEXT$9_0/m1_4800_960# TEXT$20_0/m3_9360_0# 0
C949 TEXT$22_0/m2_2880_720# TEXT$20_0/m3_2880_720# 0.23648f
C950 TEXT$21_0/m4_9360_0# TEXT$6_0/m4_7200_0# 0.03009f
C951 TEXT$21_0/m4_12960_0# TEXT$20_0/m3_12960_0# 0.40712f
C952 TEXT$1_0/m1_6000_0# TEXT$6_0/m4_4800_0# 0
C953 TEXT$4_0/m3_1200_0# TEXT$3_0/m2_1200_0# 1.11291f
C954 TEXT$23_0/m1_4320_0# TEXT$1_0/m1_2400_0# 0.00534f
C955 TEXT$21_0/m4_7920_720# TEXT$23_0/m1_7200_0# 0
C956 TEXT$23_0/m1_13680_0# TEXT$8_0/m4_9600_0# -0.00156f
C957 TEXT$22_0/m2_11700_0# TEXT$7_0/m2_6720_0# 0
C958 TEXT$4_0/m3_1200_0# TEXT$20_0/m3_4320_0# 0.0115f
C959 TEXT$1_0/m1_0_0# TEXT$3_0/m2_1200_0# 0.00488f
C960 TEXT$22_0/m2_13680_0# TEXT$22_0/m2_14400_0# 0.23093f
C961 TEXT$22_0/m2_4320_0# TEXT$22_0/m2_5760_0# 0.02095f
C962 TEXT$9_0/m1_5760_0# TEXT$20_0/m3_10080_0# 0
C963 TEXT$22_0/m2_10800_0# TEXT$23_0/m1_10800_0# 0.36457f
C964 TEXT$24_0/m3_3840_0# TEXT$9_0/m1_3840_0# 0.01435f
C965 VDD M_0/a_402461_244568# -0.01121f
C966 TEXT$23_0/m1_7920_720# TEXT$1_0/m1_4800_0# 0.00758f
C967 TEXT$21_0/m4_6480_0# TEXT$22_0/m2_5760_0# 0
C968 TEXT$1_0/m1_8400_0# TEXT$23_0/m1_10800_0# 0.02008f
C969 TEXT$21_0/m4_11700_0# TEXT$23_0/m1_11700_0# 0
C970 TEXT$24_0/m3_4800_960# TEXT$8_0/m4_4800_960# 0.42546f
C971 TEXT$1_0/m1_6000_0# TEXT$23_0/m1_8640_0# 0.01287f
C972 TEXT$23_0/m1_8640_0# TEXT$8_0/m4_3840_0# -0
C973 TEXT$21_0/m4_4320_0# TEXT$1_0/m1_2400_0# 0
C974 TEXT$23_0/m1_2160_0# TEXT$20_0/m3_2880_720# 0
C975 TEXT$8_0/m4_0_0# TEXT$22_0/m2_4320_0# 0
C976 TEXT$21_0/m4_6480_0# TEXT$21_0/m4_7200_0# 0.26312f
C977 VDD TEXT$7_0/m2_5760_0# 0.03306f
C978 TEXT$21_0/m4_6480_0# TEXT$23_0/m1_6480_0# 0
C979 TEXT$22_0/m2_7920_720# TEXT$6_0/m4_6000_0# 0
C980 TEXT$22_0/m2_4320_0# TEXT$3_0/m2_1200_0# 0.00794f
C981 TEXT$20_0/m3_2160_0# TEXT$20_0/m3_2880_720# 0.14917f
C982 TEXT$23_0/m1_10080_0# TEXT$8_0/m4_5760_0# -0.0019f
C983 TEXT$4_0/m3_10800_0# TEXT$21_0/m4_12960_0# 0
C984 TEXT$21_0/m4_17280_0# TEXT$23_0/m1_17280_0# -0
C985 TEXT$4_0/m3_9600_0# TEXT$1_0/m1_9600_0# 0.01177f
C986 TEXT$23_0/m1_7920_720# TEXT$22_0/m2_7920_720# 0.23534f
C987 TEXT$23_0/m1_9360_0# TEXT$22_0/m2_8640_0# 0.00171f
C988 TEXT$4_0/m3_9600_0# TEXT$20_0/m3_11700_0# 0.00225f
C989 TEXT$4_0/m3_6000_0# TEXT$6_0/m4_4800_0# 0.007f
C990 TEXT$1_0/m1_8400_0# TEXT$6_0/m4_9600_0# -0.00147f
C991 TEXT$1_0/m1_9600_0# TEXT$6_0/m4_8400_0# 0
C992 TEXT$6_0/m4_8400_0# TEXT$20_0/m3_11700_0# 0
C993 TEXT$8_0/m4_0_0# TEXT$7_0/m2_0_0# 0.01332f
C994 TEXT$23_0/m1_10800_0# TEXT$20_0/m3_10080_0# 0
C995 TEXT$22_0/m2_4320_0# TEXT$20_0/m3_4320_0# 0.40354f
C996 TEXT$20_0/m3_17280_0# TEXT$20_0/m3_18000_0# 0.20543f
C997 TEXT$21_0/m4_5760_0# TEXT$22_0/m2_5760_0# 0.00588f
C998 TEXT$23_0/m1_8640_0# TEXT$20_0/m3_8640_0# 0.00331f
C999 TEXT$21_0/m4_10080_0# TEXT$23_0/m1_9360_0# -0.00102f
C1000 VDD a_498947_268180# 42.48528f
C1001 TEXT$24_0/m3_4800_960# TEXT$24_0/m3_5760_0# 0.16047f
C1002 TEXT$7_0/m2_0_0# TEXT$7_0/m2_960_0# 0.16883f
C1003 TEXT$4_0/m3_4800_0# TEXT$23_0/m1_7920_720# 0
C1004 TEXT$3_0/m2_6000_0# TEXT$6_0/m4_4800_0# 0.00123f
C1005 TEXT$21_0/m4_5760_0# TEXT$23_0/m1_6480_0# -0
C1006 TEXT$23_0/m1_4320_0# TEXT$3_0/m2_2400_0# 0
C1007 TEXT$4_0/m3_8400_0# TEXT$23_0/m1_10800_0# 0
C1008 VDD TEXT$7_0/m2_4800_960# 0.00834f
C1009 TEXT$4_0/m3_2400_0# TEXT$1_0/m1_2400_0# 0.00982f
C1010 TEXT$4_0/m3_6000_0# TEXT$23_0/m1_8640_0# 0
C1011 TEXT$9_0/m1_4800_960# TEXT$8_0/m4_4800_960# 0.00249f
C1012 TEXT$24_0/m3_7680_0# TEXT$7_0/m2_7680_0# 0.7241f
C1013 TEXT$22_0/m2_15120_0# TEXT$24_0/m3_10560_0# 0
C1014 TEXT$23_0/m1_17280_0# TEXT$20_0/m3_16560_0# 0
C1015 TEXT$23_0/m1_16560_0# TEXT$20_0/m3_17280_0# 0
C1016 TEXT$6_0/m4_4800_0# TEXT$20_0/m3_7920_720# 0
C1017 TEXT$3_0/m2_0_0# TEXT$3_0/m2_1200_0# 0.20564f
C1018 TEXT$9_0/m1_9600_0# TEXT$7_0/m2_9600_0# 0.71322f
C1019 TEXT$23_0/m1_4320_0# TEXT$20_0/m3_5760_0# 0
C1020 TEXT$21_0/m4_17280_0# TEXT$21_0/m4_18000_0# 0.20695f
C1021 TEXT$7_0/m2_0_0# TEXT$20_0/m3_4320_0# 0
C1022 TEXT$23_0/m1_7920_720# TEXT$3_0/m2_4800_0# 0
C1023 TEXT$21_0/m4_5760_0# TEXT$7_0/m2_960_0# 0
C1024 TEXT$1_0/m1_1200_0# TEXT$1_0/m1_2400_0# 0.2838f
C1025 TEXT$23_0/m1_14400_0# TEXT$3_0/m2_12000_0# 0
C1026 TEXT$3_0/m2_8400_0# TEXT$23_0/m1_10800_0# 0
C1027 TEXT$3_0/m2_1200_0# TEXT$20_0/m3_3780_0# 0
C1028 TEXT$3_0/m2_6000_0# TEXT$23_0/m1_8640_0# 0
C1029 TEXT$9_0/m1_9600_0# TEXT$8_0/m4_7680_0# 0
C1030 TEXT$21_0/m4_4320_0# TEXT$3_0/m2_2400_0# 0
C1031 TEXT$23_0/m1_7920_720# TEXT$20_0/m3_7200_0# 0
C1032 TEXT$7_0/m2_2880_0# TEXT$7_0/m2_3840_0# 0.11541f
C1033 TEXT$24_0/m3_9600_0# TEXT$8_0/m4_9600_0# 0.72681f
C1034 TEXT$23_0/m1_15840_0# TEXT$23_0/m1_16560_0# 0.29377f
C1035 TEXT$20_0/m3_3780_0# TEXT$20_0/m3_4320_0# 0.13459f
C1036 TEXT$21_0/m4_4320_0# TEXT$20_0/m3_5760_0# 0
C1037 TEXT$22_0/m2_17280_0# TEXT$21_0/m4_16560_0# 0
C1038 TEXT$21_0/m4_5760_0# TEXT$20_0/m3_4320_0# 0
C1039 TEXT$1_0/m1_4800_0# TEXT$23_0/m1_7200_0# 0.01631f
C1040 TEXT$21_0/m4_10080_0# TEXT$23_0/m1_10080_0# -0
C1041 TEXT$24_0/m3_0_0# VDD 0.00863f
C1042 TEXT$7_0/m2_10560_0# TEXT$20_0/m3_14400_0# 0.0016f
C1043 TEXT$4_0/m3_8400_0# TEXT$6_0/m4_9600_0# 0.00209f
C1044 TEXT$4_0/m3_9600_0# TEXT$6_0/m4_8400_0# 0.00894f
C1045 TEXT$22_0/m2_15840_0# TEXT$20_0/m3_16560_0# 0.00184f
C1046 TEXT$24_0/m3_5760_0# TEXT$9_0/m1_4800_960# 0
C1047 TEXT$21_0/m4_11700_0# TEXT$24_0/m3_6720_0# 0
C1048 TEXT$7_0/m2_2880_0# TEXT$8_0/m4_2160_0# 0
C1049 TEXT$3_0/m2_8400_0# TEXT$6_0/m4_9600_0# 0
C1050 TEXT$9_0/m1_6720_0# TEXT$20_0/m3_11700_0# 0
C1051 TEXT$6_0/m4_0_0# TEXT$23_0/m1_2880_720# 0
C1052 TEXT$23_0/m1_13680_0# TEXT$7_0/m2_9600_0# 0.00219f
C1053 TEXT$22_0/m2_15120_0# TEXT$23_0/m1_15840_0# 0.00132f
C1054 TEXT$21_0/m4_6480_0# TEXT$1_0/m1_3600_0# 0
C1055 TEXT$8_0/m4_10560_0# TEXT$8_0/m4_9600_0# 0.17706f
C1056 TEXT$22_0/m2_9360_0# TEXT$6_0/m4_7200_0# 0
C1057 TEXT$22_0/m2_7920_720# TEXT$23_0/m1_7200_0# 0
C1058 TEXT$1_0/m1_10800_0# TEXT$20_0/m3_12960_0# 0
C1059 TEXT$21_0/m4_13680_0# TEXT$20_0/m3_13680_0# 0.34758f
C1060 TEXT$1_0/m1_7200_0# TEXT$6_0/m4_6000_0# 0
C1061 TEXT$4_0/m3_2400_0# TEXT$3_0/m2_2400_0# 1.00682f
C1062 TEXT$21_0/m4_720_0# TEXT$20_0/m3_0_0# 0
C1063 TEXT$7_0/m2_2160_0# TEXT$7_0/m2_2880_0# 0.10378f
C1064 TEXT$24_0/m3_0_0# TEXT$22_0/m2_4320_0# 0
C1065 TEXT$1_0/m1_1200_0# TEXT$3_0/m2_2400_0# 0.007f
C1066 TEXT$22_0/m2_5760_0# TEXT$22_0/m2_6480_0# 0.15515f
C1067 TEXT$22_0/m2_14400_0# TEXT$22_0/m2_15120_0# 0.2155f
C1068 TEXT$4_0/m3_4800_0# TEXT$23_0/m1_7200_0# 0
C1069 TEXT$24_0/m3_4800_960# TEXT$9_0/m1_4800_960# 0.00768f
C1070 TEXT$23_0/m1_6480_0# TEXT$8_0/m4_2160_0# 0
C1071 TEXT$21_0/m4_7200_0# TEXT$22_0/m2_6480_0# 0
C1072 TEXT$22_0/m2_11700_0# TEXT$8_0/m4_7680_0# 0
C1073 TEXT$1_0/m1_2400_0# TEXT$20_0/m3_4320_0# 0
C1074 TEXT$1_0/m1_9600_0# TEXT$23_0/m1_11700_0# 0.00115f
C1075 TEXT$21_0/m4_12960_0# TEXT$23_0/m1_12960_0# -0
C1076 TEXT$23_0/m1_6480_0# TEXT$22_0/m2_6480_0# 0.40242f
C1077 TEXT$23_0/m1_11700_0# TEXT$20_0/m3_11700_0# 0.00157f
C1078 TEXT$21_0/m4_5760_0# TEXT$1_0/m1_3600_0# -0
C1079 TEXT$3_0/m2_4800_0# TEXT$23_0/m1_7200_0# 0
C1080 TEXT$21_0/m4_7200_0# TEXT$21_0/m4_7920_720# 0.12576f
C1081 TEXT$7_0/m2_960_0# TEXT$8_0/m4_2160_0# 0
C1082 VDD TEXT$7_0/m2_7680_0# 0.01668f
C1083 TEXT$22_0/m2_13680_0# TEXT$8_0/m4_9600_0# 0
C1084 TEXT$23_0/m1_5760_0# TEXT$6_0/m4_3600_0# -0
C1085 TEXT$9_0/m1_0_0# VDD 0.03274f
C1086 TEXT$4_0/m3_3600_0# TEXT$21_0/m4_6480_0# 0
C1087 TEXT$24_0/m3_0_0# TEXT$7_0/m2_0_0# 0.59794f
C1088 TEXT$20_0/m3_7200_0# TEXT$23_0/m1_7200_0# 0.00299f
C1089 TEXT$22_0/m2_11700_0# TEXT$21_0/m4_11700_0# 0.00207f
C1090 TEXT$4_0/m3_10800_0# TEXT$1_0/m1_10800_0# 0.01242f
C1091 TEXT$23_0/m1_6480_0# TEXT$7_0/m2_2160_0# 0
C1092 TEXT$23_0/m1_9360_0# TEXT$22_0/m2_10080_0# 0
C1093 TEXT$4_0/m3_10800_0# TEXT$20_0/m3_12960_0# 0.0125f
C1094 TEXT$4_0/m3_7200_0# TEXT$6_0/m4_6000_0# 0.00978f
C1095 TEXT$1_0/m1_10800_0# TEXT$6_0/m4_9600_0# 0
C1096 TEXT$1_0/m1_9600_0# TEXT$6_0/m4_10800_0# 0
C1097 TEXT$21_0/m4_6480_0# TEXT$3_0/m2_3600_0# 0
C1098 TEXT$22_0/m2_5760_0# TEXT$20_0/m3_5760_0# 0.41032f
C1099 TEXT$23_0/m1_9360_0# TEXT$1_0/m1_7200_0# 0.01782f
C1100 TEXT$21_0/m4_6480_0# TEXT$20_0/m3_6480_0# 0.40538f
C1101 TEXT$7_0/m2_960_0# TEXT$7_0/m2_2160_0# 0.10378f
C1102 TEXT$23_0/m1_6480_0# TEXT$20_0/m3_5760_0# 0
C1103 TEXT$3_0/m2_7200_0# TEXT$6_0/m4_6000_0# 0.0019f
C1104 TEXT$8_0/m4_3840_0# VDD 0.00998f
C1105 TEXT$24_0/m3_3840_0# TEXT$23_0/m1_8640_0# 0
C1106 TEXT$22_0/m2_17280_0# TEXT$21_0/m4_17280_0# 0.00593f
C1107 TEXT$4_0/m3_3600_0# TEXT$21_0/m4_5760_0# 0
C1108 TEXT$23_0/m1_11700_0# TEXT$6_0/m4_8400_0# 0
C1109 TEXT$3_0/m2_9600_0# TEXT$3_0/m2_10800_0# 0.12477f
C1110 TEXT$24_0/m3_9600_0# TEXT$7_0/m2_9600_0# 0.71411f
C1111 TEXT$23_0/m1_18000_0# TEXT$20_0/m3_17280_0# 0
C1112 TEXT$3_0/m2_1200_0# TEXT$3_0/m2_2400_0# 0.25104f
C1113 TEXT$9_0/m1_10560_0# TEXT$7_0/m2_10560_0# 0.74016f
C1114 TEXT$7_0/m2_960_0# TEXT$20_0/m3_5760_0# 0
C1115 TEXT$21_0/m4_8640_0# TEXT$21_0/m4_9360_0# 0.26312f
C1116 TEXT$22_0/m2_4320_0# TEXT$9_0/m1_0_0# 0
C1117 TEXT$1_0/m1_2400_0# TEXT$1_0/m1_3600_0# 0.21322f
C1118 TEXT$24_0/m3_9600_0# TEXT$8_0/m4_7680_0# 0
C1119 TEXT$21_0/m4_8640_0# TEXT$7_0/m2_4800_960# 0
C1120 TEXT$3_0/m2_2400_0# TEXT$20_0/m3_4320_0# 0
C1121 TEXT$21_0/m4_5760_0# TEXT$3_0/m2_3600_0# 0
C1122 VDD a_499016_248165# 41.80168f
C1123 TEXT$23_0/m1_10080_0# TEXT$22_0/m2_10080_0# 0.40191f
C1124 TEXT$23_0/m1_9360_0# TEXT$20_0/m3_9360_0# 0.00288f
C1125 TEXT$7_0/m2_3840_0# TEXT$7_0/m2_4800_960# 0.11044f
C1126 TEXT$23_0/m1_16560_0# TEXT$23_0/m1_17280_0# 0.1367f
C1127 TEXT$20_0/m3_4320_0# TEXT$20_0/m3_5760_0# 0.03005f
C1128 TEXT$21_0/m4_5760_0# TEXT$20_0/m3_6480_0# 0
C1129 TEXT$23_0/m1_10080_0# TEXT$1_0/m1_7200_0# 0.01234f
C1130 TEXT$24_0/m3_2160_0# VDD 0.00368f
C1131 TEXT$4_0/m3_9600_0# TEXT$6_0/m4_10800_0# 0
C1132 TEXT$4_0/m3_10800_0# TEXT$6_0/m4_9600_0# 0.00318f
C1133 TEXT$22_0/m2_17280_0# TEXT$20_0/m3_16560_0# 0
C1134 TEXT$22_0/m2_16560_0# TEXT$20_0/m3_17280_0# 0.00101f
C1135 TEXT$8_0/m4_10560_0# TEXT$7_0/m2_9600_0# 0.0011f
C1136 TEXT$21_0/m4_18000_0# TEXT$20_0/m3_18000_0# 0.34763f
C1137 TEXT$9_0/m1_0_0# TEXT$7_0/m2_0_0# 0.59211f
C1138 TEXT$22_0/m2_14400_0# TEXT$3_0/m2_12000_0# 0.02147f
C1139 TEXT$24_0/m3_6720_0# TEXT$20_0/m3_11700_0# 0.00136f
C1140 TEXT$9_0/m1_7680_0# TEXT$8_0/m4_6720_0# -0
C1141 TEXT$21_0/m4_13680_0# TEXT$9_0/m1_9600_0# 0
C1142 TEXT$22_0/m2_6480_0# TEXT$1_0/m1_3600_0# 0
C1143 TEXT$23_0/m1_14400_0# TEXT$7_0/m2_10560_0# 0.0021f
C1144 TEXT$24_0/m3_5760_0# TEXT$24_0/m3_6720_0# 0.21746f
C1145 TEXT$21_0/m4_7200_0# TEXT$1_0/m1_4800_0# 0
C1146 TEXT$23_0/m1_9360_0# TEXT$3_0/m2_7200_0# 0
C1147 TEXT$22_0/m2_15840_0# TEXT$23_0/m1_16560_0# 0.00171f
C1148 TEXT$9_0/m1_3840_0# TEXT$23_0/m1_8640_0# 0.00868f
C1149 TEXT$8_0/m4_5760_0# TEXT$7_0/m2_5760_0# 0.01366f
C1150 TEXT$23_0/m1_10080_0# TEXT$20_0/m3_9360_0# 0
C1151 TEXT$4_0/m3_3600_0# TEXT$1_0/m1_2400_0# 0.00143f
C1152 TEXT$21_0/m4_15120_0# TEXT$1_0/m1_12000_0# -0
C1153 TEXT$21_0/m4_14400_0# TEXT$20_0/m3_14400_0# 0.40882f
C1154 TEXT$1_0/m1_8400_0# TEXT$6_0/m4_7200_0# 0
C1155 TEXT$23_0/m1_11700_0# TEXT$9_0/m1_6720_0# 0.00106f
C1156 TEXT$20_0/m3_0_0# TEXT$20_0/m3_720_0# 0.2313f
C1157 TEXT$7_0/m2_5760_0# TEXT$7_0/m2_6720_0# 0.17804f
C1158 TEXT$24_0/m3_960_0# TEXT$22_0/m2_5760_0# 0
C1159 TEXT$22_0/m2_13680_0# TEXT$7_0/m2_9600_0# 0.01326f
C1160 TEXT$1_0/m1_2400_0# TEXT$3_0/m2_3600_0# 0.00446f
C1161 TEXT$22_0/m2_15120_0# TEXT$22_0/m2_15840_0# 0.18145f
C1162 TEXT$22_0/m2_6480_0# TEXT$22_0/m2_7200_0# 0.22232f
C1163 TEXT$24_0/m3_2880_0# TEXT$23_0/m1_7200_0# 0
C1164 TEXT$21_0/m4_0_0# TEXT$22_0/m2_0_0# 0.00474f
C1165 TEXT$21_0/m4_7920_720# TEXT$22_0/m2_7200_0# 0
C1166 TEXT$21_0/m4_6480_0# TEXT$24_0/m3_2160_0# 0
C1167 TEXT$21_0/m4_13680_0# TEXT$23_0/m1_13680_0# 0
C1168 TEXT$1_0/m1_10800_0# TEXT$23_0/m1_12960_0# 0.00794f
C1169 TEXT$22_0/m2_2160_0# TEXT$6_0/m4_0_0# 0
C1170 TEXT$23_0/m1_12960_0# TEXT$20_0/m3_12960_0# 0.00329f
C1171 TEXT$20_0/m3_7200_0# TEXT$7_0/m2_2880_0# 0.00101f
C1172 TEXT$4_0/m3_3600_0# TEXT$22_0/m2_6480_0# 0
C1173 TEXT$23_0/m1_10080_0# TEXT$3_0/m2_7200_0# 0
C1174 TEXT$8_0/m4_0_0# TEXT$24_0/m3_960_0# 0.0052f
C1175 VDD TEXT$7_0/m2_10560_0# 0.02937f
C1176 TEXT$23_0/m1_9360_0# TEXT$8_0/m4_4800_960# -0
C1177 TEXT$8_0/m4_5760_0# TEXT$7_0/m2_4800_960# 0
C1178 TEXT$9_0/m1_2160_0# VDD 0.01552f
C1179 TEXT$6_0/m4_7200_0# TEXT$20_0/m3_10080_0# 0
C1180 PU PD 0.34623f
C1181 TEXT$4_0/m3_4800_0# TEXT$21_0/m4_7200_0# 0
C1182 TEXT$24_0/m3_960_0# TEXT$7_0/m2_960_0# 0.65629f
C1183 TEXT$22_0/m2_6480_0# TEXT$3_0/m2_3600_0# 0.01056f
C1184 TEXT$21_0/m4_10080_0# TEXT$7_0/m2_5760_0# 0
C1185 TEXT$20_0/m3_6480_0# TEXT$8_0/m4_2160_0# 0
C1186 TEXT$22_0/m2_11700_0# TEXT$1_0/m1_9600_0# 0
C1187 TEXT$22_0/m2_12960_0# TEXT$21_0/m4_12960_0# 0.00591f
C1188 TEXT$4_0/m3_12000_0# TEXT$21_0/m4_15120_0# 0
C1189 TEXT$4_0/m3_12000_0# TEXT$1_0/m1_12000_0# 0.01556f
C1190 TEXT$22_0/m2_11700_0# TEXT$20_0/m3_11700_0# 0.1943f
C1191 TEXT$21_0/m4_14400_0# TEXT$6_0/m4_12000_0# 0.03241f
C1192 TEXT$4_0/m3_8400_0# TEXT$6_0/m4_7200_0# 0.00184f
C1193 TEXT$1_0/m1_10800_0# TEXT$6_0/m4_12000_0# -0.00146f
C1194 TEXT$1_0/m1_12000_0# TEXT$6_0/m4_10800_0# 0
C1195 TEXT$21_0/m4_7200_0# TEXT$3_0/m2_4800_0# 0
C1196 TEXT$22_0/m2_6480_0# TEXT$20_0/m3_6480_0# 0.40709f
C1197 TEXT$21_0/m4_5760_0# TEXT$24_0/m3_2160_0# 0
C1198 TEXT$23_0/m1_2880_720# TEXT$23_0/m1_3780_0# 0.06713f
C1199 TEXT$21_0/m4_7200_0# TEXT$20_0/m3_7200_0# 0.36636f
C1200 TEXT$9_0/m1_2880_0# TEXT$23_0/m1_7200_0# 0.02195f
C1201 TEXT$24_0/m3_5760_0# TEXT$23_0/m1_9360_0# 0
C1202 TEXT$21_0/m4_2880_720# TEXT$6_0/m4_0_0# 0.01349f
C1203 TEXT$3_0/m2_8400_0# TEXT$6_0/m4_7200_0# 0
C1204 TEXT$4_0/m3_3600_0# TEXT$20_0/m3_5760_0# 0.016f
C1205 TEXT$21_0/m4_9360_0# TEXT$22_0/m2_8640_0# 0
C1206 TEXT$3_0/m2_10800_0# TEXT$3_0/m2_12000_0# 0.11662f
C1207 TEXT$8_0/m4_2880_0# VDD 0.00729f
C1208 TEXT$24_0/m3_10560_0# TEXT$7_0/m2_10560_0# 0.74066f
C1209 TEXT$4_0/m3_1200_0# TEXT$6_0/m4_0_0# 0.007f
C1210 TEXT$3_0/m2_2400_0# TEXT$3_0/m2_3600_0# 0.18694f
C1211 TEXT$22_0/m2_8640_0# TEXT$7_0/m2_4800_960# 0.01072f
C1212 TEXT$7_0/m2_2160_0# TEXT$20_0/m3_6480_0# 0
C1213 TEXT$21_0/m4_8640_0# TEXT$1_0/m1_6000_0# -0
C1214 TEXT$1_0/m1_3600_0# TEXT$1_0/m1_4800_0# 0.29851f
C1215 TEXT$21_0/m4_9360_0# TEXT$21_0/m4_10080_0# 0.11931f
C1216 TEXT$21_0/m4_8640_0# TEXT$8_0/m4_3840_0# 0.00737f
C1217 TEXT$1_0/m1_0_0# TEXT$6_0/m4_0_0# 0.00594f
C1218 TEXT$3_0/m2_3600_0# TEXT$20_0/m3_5760_0# 0
C1219 TEXT$8_0/m4_3840_0# TEXT$7_0/m2_3840_0# 0.01633f
C1220 TEXT$21_0/m4_6480_0# TEXT$9_0/m1_2160_0# 0
C1221 TEXT$24_0/m3_6720_0# TEXT$9_0/m1_6720_0# 0.01099f
C1222 TEXT$21_0/m4_10800_0# TEXT$20_0/m3_10800_0# 0.36602f
C1223 TEXT$22_0/m2_11700_0# TEXT$4_0/m3_9600_0# 0
C1224 TEXT$23_0/m1_17280_0# TEXT$23_0/m1_18000_0# 0.22968f
C1225 TEXT$20_0/m3_5760_0# TEXT$20_0/m3_6480_0# 0.18616f
C1226 TEXT$22_0/m2_11700_0# TEXT$6_0/m4_8400_0# 0
C1227 TEXT$8_0/m4_0_0# TEXT$9_0/m1_960_0# -0
C1228 TEXT$22_0/m2_18000_0# TEXT$20_0/m3_17280_0# 0
C1229 TEXT$22_0/m2_17280_0# TEXT$20_0/m3_18000_0# 0.00261f
C1230 TEXT$4_0/m3_10800_0# TEXT$6_0/m4_12000_0# 0
C1231 TEXT$4_0/m3_12000_0# TEXT$6_0/m4_10800_0# 0.00415f
C1232 TEXT$9_0/m1_960_0# TEXT$7_0/m2_960_0# 0.65326f
C1233 TEXT$24_0/m3_4800_960# TEXT$23_0/m1_9360_0# 0
C1234 TEXT$24_0/m3_5760_0# TEXT$23_0/m1_10080_0# 0
C1235 TEXT$24_0/m3_7680_0# TEXT$8_0/m4_6720_0# 0.00734f
C1236 TEXT$21_0/m4_13680_0# TEXT$24_0/m3_9600_0# 0
C1237 TEXT$21_0/m4_14400_0# TEXT$9_0/m1_10560_0# 0
C1238 TEXT$22_0/m2_7200_0# TEXT$1_0/m1_4800_0# 0
C1239 TEXT$21_0/m4_8640_0# TEXT$20_0/m3_8640_0# 0.40548f
C1240 TEXT$24_0/m3_3840_0# VDD 0.00687f
C1241 TEXT$9_0/m1_9600_0# TEXT$20_0/m3_13680_0# 0
C1242 TEXT$22_0/m2_3780_0# TEXT$6_0/m4_1200_0# 0
C1243 TEXT$20_0/m3_8640_0# TEXT$7_0/m2_3840_0# 0
C1244 TEXT$22_0/m2_17280_0# TEXT$23_0/m1_16560_0# 0
C1245 TEXT$22_0/m2_16560_0# TEXT$23_0/m1_17280_0# 0
C1246 TEXT$21_0/m4_7920_720# TEXT$8_0/m4_3840_0# 0.01068f
C1247 TEXT$21_0/m4_18000_0# TEXT$23_0/m1_18000_0# 0
C1248 TEXT$4_0/m3_6000_0# TEXT$21_0/m4_8640_0# 0
C1249 TEXT$4_0/m3_4800_0# TEXT$1_0/m1_3600_0# 0.00256f
C1250 TEXT$24_0/m3_6720_0# TEXT$23_0/m1_11700_0# 0
C1251 TEXT$1_0/m1_12000_0# TEXT$20_0/m3_15120_0# 0
C1252 TEXT$21_0/m4_15120_0# TEXT$20_0/m3_15120_0# 0.36602f
C1253 TEXT$24_0/m3_2880_0# TEXT$7_0/m2_2880_0# 0.65407f
C1254 TEXT$24_0/m3_2160_0# TEXT$8_0/m4_2160_0# 0.3512f
C1255 TEXT$23_0/m1_4320_0# TEXT$6_0/m4_1200_0# 0
C1256 TEXT$21_0/m4_11700_0# TEXT$3_0/m2_9600_0# 0
C1257 TEXT$7_0/m2_6720_0# TEXT$7_0/m2_7680_0# 0.24926f
C1258 TEXT$24_0/m3_2160_0# TEXT$22_0/m2_6480_0# 0
C1259 TEXT$22_0/m2_14400_0# TEXT$7_0/m2_10560_0# 0.00732f
C1260 TEXT$1_0/m1_3600_0# TEXT$3_0/m2_4800_0# 0.00675f
C1261 TEXT$21_0/m4_8640_0# TEXT$3_0/m2_6000_0# 0
C1262 TEXT$22_0/m2_7200_0# TEXT$22_0/m2_7920_720# 0.09293f
C1263 TEXT$22_0/m2_15840_0# TEXT$22_0/m2_16560_0# 0.22232f
C1264 TEXT$3_0/m2_0_0# TEXT$6_0/m4_0_0# 0.0087f
C1265 TEXT$24_0/m3_0_0# TEXT$24_0/m3_960_0# 0.21166f
C1266 TEXT$21_0/m4_720_0# TEXT$22_0/m2_720_0# 0.00321f
C1267 TEXT$21_0/m4_8640_0# TEXT$20_0/m3_7920_720# 0
C1268 TEXT$21_0/m4_14400_0# TEXT$23_0/m1_14400_0# -0
C1269 TEXT$23_0/m1_13680_0# TEXT$20_0/m3_13680_0# 0.00233f
C1270 TEXT$23_0/m1_9360_0# TEXT$9_0/m1_4800_960# 0.00982f
C1271 TEXT$20_0/m3_7920_720# TEXT$7_0/m2_3840_0# 0
C1272 TEXT$22_0/m2_11700_0# TEXT$9_0/m1_6720_0# 0
C1273 TEXT$21_0/m4_4320_0# TEXT$6_0/m4_1200_0# 0.01309f
C1274 TEXT$4_0/m3_4800_0# TEXT$22_0/m2_7200_0# 0
C1275 TEXT$8_0/m4_9600_0# TEXT$7_0/m2_7680_0# 0
C1276 TEXT$9_0/m1_3840_0# VDD 0.0314f
C1277 TEXT$23_0/m1_4320_0# TEXT$23_0/m1_5760_0# 0.01943f
C1278 TEXT$4_0/m3_6000_0# TEXT$21_0/m4_7920_720# 0
C1279 TEXT$24_0/m3_2160_0# TEXT$7_0/m2_2160_0# 0.34994f
C1280 TEXT$24_0/m3_2880_0# TEXT$21_0/m4_7200_0# 0
C1281 TEXT$22_0/m2_10080_0# TEXT$7_0/m2_5760_0# 0.01611f
C1282 TEXT$24_0/m3_2880_0# TEXT$23_0/m1_6480_0# 0
C1283 TEXT$21_0/m4_0_0# TEXT$23_0/m1_0_0# -0
C1284 TEXT$22_0/m2_7200_0# TEXT$3_0/m2_4800_0# 0.01754f
C1285 VDD VIN 19.90989f
C1286 TEXT$21_0/m4_10800_0# TEXT$7_0/m2_6720_0# 0
C1287 TEXT$4_0/m3_3600_0# TEXT$4_0/m3_4800_0# 0.32982f
C1288 TEXT$9_0/m1_5760_0# VDD 0.03045f
C1289 TEXT$22_0/m2_12960_0# TEXT$1_0/m1_10800_0# 0
C1290 TEXT$22_0/m2_13680_0# TEXT$21_0/m4_13680_0# 0.00319f
C1291 TEXT$22_0/m2_12960_0# TEXT$20_0/m3_12960_0# 0.41002f
C1292 TEXT$4_0/m3_12000_0# TEXT$20_0/m3_15120_0# 0.01053f
C1293 TEXT$21_0/m4_7920_720# TEXT$3_0/m2_6000_0# 0
C1294 TEXT$22_0/m2_7200_0# TEXT$20_0/m3_7200_0# 0.36732f
C1295 TEXT$6_0/m4_12000_0# TEXT$20_0/m3_14400_0# 0
C1296 TEXT$9_0/m1_2880_0# TEXT$7_0/m2_2880_0# 0.65157f
C1297 TEXT$21_0/m4_4320_0# TEXT$23_0/m1_5760_0# -0
C1298 TEXT$24_0/m3_2160_0# TEXT$20_0/m3_5760_0# 0
C1299 TEXT$21_0/m4_7920_720# TEXT$20_0/m3_7920_720# 0.23623f
C1300 TEXT$6_0/m4_0_0# TEXT$20_0/m3_2880_720# 0
C1301 TEXT$22_0/m2_8640_0# TEXT$22_0/m2_9360_0# 0.22232f
C1302 TEXT$22_0/m2_0_0# TEXT$23_0/m1_0_0# 0.44019f
C1303 TEXT$8_0/m4_6720_0# VDD 0.01061f
C1304 TEXT$22_0/m2_11700_0# TEXT$23_0/m1_11700_0# 0.19314f
C1305 TEXT$21_0/m4_9360_0# TEXT$22_0/m2_10080_0# 0
C1306 TEXT$21_0/m4_10080_0# TEXT$22_0/m2_9360_0# 0
C1307 TEXT$4_0/m3_1200_0# TEXT$6_0/m4_2400_0# 0.0323f
C1308 TEXT$4_0/m3_2400_0# TEXT$6_0/m4_1200_0# 0.00978f
C1309 TEXT$22_0/m2_8640_0# TEXT$1_0/m1_6000_0# 0
C1310 TEXT$9_0/m1_2160_0# TEXT$8_0/m4_2160_0# 0.00147f
C1311 TEXT$22_0/m2_8640_0# TEXT$8_0/m4_3840_0# 0
C1312 TEXT$3_0/m2_3600_0# TEXT$3_0/m2_4800_0# 0.26172f
C1313 TEXT$22_0/m2_6480_0# TEXT$9_0/m1_2160_0# 0
C1314 TEXT$21_0/m4_9360_0# TEXT$1_0/m1_7200_0# -0
C1315 TEXT$1_0/m1_4800_0# TEXT$1_0/m1_6000_0# 0.23454f
C1316 TEXT$21_0/m4_10080_0# TEXT$21_0/m4_10800_0# 0.24565f
C1317 VDD VCM_OUT 0.12526f
C1318 TEXT$24_0/m3_960_0# TEXT$9_0/m1_0_0# 0
C1319 TEXT$24_0/m3_0_0# TEXT$9_0/m1_960_0# 0
C1320 TEXT$1_0/m1_1200_0# TEXT$6_0/m4_1200_0# 0.00486f
C1321 TEXT$22_0/m2_10800_0# TEXT$20_0/m3_10800_0# 0.36742f
C1322 TEXT$24_0/m3_7680_0# TEXT$9_0/m1_7680_0# 0.00861f
C1323 TEXT$21_0/m4_7200_0# TEXT$9_0/m1_2880_0# -0
C1324 TEXT$8_0/m4_2880_0# TEXT$7_0/m2_3840_0# 0
C1325 TEXT$22_0/m2_12960_0# TEXT$4_0/m3_10800_0# 0
C1326 TEXT$20_0/m3_6480_0# TEXT$20_0/m3_7200_0# 0.26159f
C1327 TEXT$21_0/m4_3780_0# TEXT$23_0/m1_3780_0# 0
C1328 TEXT$9_0/m1_2160_0# TEXT$7_0/m2_2160_0# 0.34642f
C1329 TEXT$22_0/m2_8640_0# TEXT$20_0/m3_8640_0# 0.40628f
C1330 TEXT$21_0/m4_14400_0# TEXT$24_0/m3_10560_0# 0
C1331 TEXT$22_0/m2_1440_0# TEXT$22_0/m2_720_0# 0.23093f
C1332 TEXT$24_0/m3_9600_0# TEXT$20_0/m3_13680_0# 0.02434f
C1333 TEXT$22_0/m2_7920_720# TEXT$8_0/m4_3840_0# 0
C1334 TEXT$21_0/m4_9360_0# TEXT$20_0/m3_9360_0# 0.42035f
C1335 TEXT$22_0/m2_7920_720# TEXT$1_0/m1_6000_0# 0
C1336 TEXT$9_0/m1_10560_0# TEXT$20_0/m3_14400_0# 0
C1337 TEXT$22_0/m2_4320_0# TEXT$6_0/m4_2400_0# 0
C1338 TEXT$8_0/m4_2880_0# TEXT$8_0/m4_2160_0# 0.15081f
C1339 TEXT$20_0/m3_9360_0# TEXT$7_0/m2_4800_960# 0
C1340 TEXT$22_0/m2_18000_0# TEXT$23_0/m1_17280_0# 0
C1341 TEXT$22_0/m2_17280_0# TEXT$23_0/m1_18000_0# 0.00175f
C1342 TEXT$4_0/m3_6000_0# TEXT$22_0/m2_8640_0# 0
C1343 TEXT$21_0/m4_720_0# TEXT$20_0/m3_720_0# 0.34763f
C1344 TEXT$4_0/m3_7200_0# TEXT$21_0/m4_9360_0# 0
C1345 TEXT$4_0/m3_6000_0# TEXT$1_0/m1_4800_0# 0.00156f
C1346 TEXT$20_0/m3_10080_0# TEXT$20_0/m3_10800_0# 0.24398f
C1347 TEXT$24_0/m3_3840_0# TEXT$21_0/m4_8640_0# 0.00225f
C1348 TEXT$21_0/m4_15840_0# TEXT$20_0/m3_15840_0# 0.40604f
C1349 TEXT$24_0/m3_3840_0# TEXT$7_0/m2_3840_0# 0.72679f
C1350 TEXT$23_0/m1_13680_0# TEXT$9_0/m1_9600_0# 0.0153f
C1351 TEXT$22_0/m2_2160_0# TEXT$23_0/m1_2880_720# 0
C1352 TEXT$22_0/m2_8640_0# TEXT$3_0/m2_6000_0# 0.01379f
C1353 TEXT$21_0/m4_15120_0# TEXT$8_0/m4_10560_0# 0.02842f
C1354 TEXT$21_0/m4_3780_0# TEXT$23_0/m1_2880_720# 0
C1355 TEXT$23_0/m1_5760_0# TEXT$22_0/m2_5760_0# 0.40253f
C1356 TEXT$4_0/m3_8400_0# TEXT$20_0/m3_10800_0# 0.03206f
C1357 TEXT$21_0/m4_12960_0# TEXT$3_0/m2_10800_0# 0
C1358 TEXT$1_0/m1_9600_0# TEXT$3_0/m2_9600_0# 1.01481f
C1359 TEXT$7_0/m2_7680_0# TEXT$7_0/m2_9600_0# 0.02237f
C1360 TEXT$21_0/m4_9360_0# TEXT$3_0/m2_7200_0# 0
C1361 TEXT$20_0/m3_11700_0# TEXT$3_0/m2_9600_0# 0
C1362 TEXT$1_0/m1_4800_0# TEXT$3_0/m2_6000_0# 0.00488f
C1363 TEXT$22_0/m2_16560_0# TEXT$22_0/m2_17280_0# 0.10328f
C1364 TEXT$7_0/m2_2160_0# TEXT$8_0/m4_2880_0# 0
C1365 TEXT$22_0/m2_7920_720# TEXT$20_0/m3_8640_0# 0
C1366 TEXT$4_0/m3_1200_0# TEXT$23_0/m1_3780_0# 0
C1367 TEXT$3_0/m2_1200_0# TEXT$6_0/m4_1200_0# 0.0097f
C1368 TEXT$24_0/m3_960_0# TEXT$24_0/m3_2160_0# 0.14271f
C1369 TEXT$22_0/m2_720_0# TEXT$20_0/m3_720_0# 0.34869f
C1370 TEXT$22_0/m2_18000_0# TEXT$21_0/m4_18000_0# 0.00321f
C1371 TEXT$9_0/m1_0_0# TEXT$9_0/m1_960_0# 0.19747f
C1372 TEXT$23_0/m1_7920_720# TEXT$6_0/m4_6000_0# 0
C1373 TEXT$8_0/m4_4800_960# TEXT$7_0/m2_5760_0# 0
C1374 TEXT$8_0/m4_7680_0# TEXT$7_0/m2_7680_0# 0.01302f
C1375 TEXT$1_0/m1_4800_0# TEXT$20_0/m3_7920_720# 0
C1376 TEXT$1_0/m1_12000_0# TEXT$23_0/m1_15120_0# 0.00684f
C1377 TEXT$21_0/m4_15120_0# TEXT$23_0/m1_15120_0# 0
C1378 TEXT$23_0/m1_6480_0# TEXT$23_0/m1_5760_0# 0.20758f
C1379 TEXT$22_0/m2_11700_0# TEXT$24_0/m3_6720_0# 0
C1380 TEXT$6_0/m4_1200_0# TEXT$20_0/m3_4320_0# 0
C1381 TEXT$23_0/m1_14400_0# TEXT$20_0/m3_14400_0# 0.00303f
C1382 TEXT$3_0/m2_8400_0# TEXT$20_0/m3_10800_0# 0
C1383 TEXT$24_0/m3_2880_0# TEXT$22_0/m2_7200_0# 0
C1384 TEXT$4_0/m3_6000_0# TEXT$22_0/m2_7920_720# 0
C1385 TEXT$21_0/m4_720_0# TEXT$23_0/m1_720_0# 0
C1386 TEXT$8_0/m4_9600_0# TEXT$7_0/m2_10560_0# 0
C1387 TEXT$8_0/m4_0_0# TEXT$8_0/m4_960_0# 0.21726f
C1388 TEXT$23_0/m1_5760_0# TEXT$7_0/m2_960_0# 0
C1389 TEXT$22_0/m2_10800_0# TEXT$7_0/m2_6720_0# 0.01349f
C1390 TEXT$24_0/m3_3840_0# TEXT$21_0/m4_7920_720# 0
C1391 TEXT$8_0/m4_960_0# TEXT$7_0/m2_960_0# 0.01366f
C1392 TEXT$22_0/m2_7920_720# TEXT$3_0/m2_6000_0# 0.00926f
C1393 TEXT$4_0/m3_4800_0# TEXT$4_0/m3_6000_0# 0.25914f
C1394 TEXT$9_0/m1_7680_0# VDD 0.01562f
C1395 TEXT$21_0/m4_2880_720# TEXT$23_0/m1_2880_720# 0
C1396 TEXT$22_0/m2_14400_0# TEXT$21_0/m4_14400_0# 0.00431f
C1397 TEXT$21_0/m4_8640_0# TEXT$9_0/m1_3840_0# -0.00427f
C1398 TEXT$22_0/m2_13680_0# TEXT$20_0/m3_13680_0# 0.34869f
C1399 TEXT$23_0/m1_5760_0# TEXT$20_0/m3_4320_0# 0
C1400 TEXT$22_0/m2_7920_720# TEXT$20_0/m3_7920_720# 0.23648f
C1401 TEXT$9_0/m1_3840_0# TEXT$7_0/m2_3840_0# 0.72194f
C1402 TEXT$24_0/m3_5760_0# TEXT$7_0/m2_5760_0# 0.65629f
C1403 TEXT$23_0/m1_720_0# TEXT$22_0/m2_720_0# 0.34645f
C1404 TEXT$21_0/m4_9360_0# TEXT$8_0/m4_4800_960# 0.02245f
C1405 TEXT$22_0/m2_4320_0# TEXT$23_0/m1_3780_0# 0
C1406 TEXT$4_0/m3_9600_0# TEXT$3_0/m2_9600_0# 1.00825f
C1407 TEXT$8_0/m4_4800_960# TEXT$7_0/m2_4800_960# 0.00883f
C1408 TEXT$6_0/m4_8400_0# TEXT$3_0/m2_9600_0# 0.00205f
C1409 TEXT$8_0/m4_5760_0# TEXT$20_0/m3_10080_0# 0.00139f
C1410 TEXT$1_0/m1_0_0# TEXT$23_0/m1_2880_720# 0.00794f
C1411 TEXT$22_0/m2_9360_0# TEXT$22_0/m2_10080_0# 0.10113f
C1412 TEXT$4_0/m3_4800_0# TEXT$20_0/m3_7920_720# 0.0115f
C1413 TEXT$22_0/m2_12960_0# TEXT$23_0/m1_12960_0# 0.40251f
C1414 TEXT$4_0/m3_12000_0# TEXT$23_0/m1_15120_0# 0
C1415 TEXT$24_0/m3_2880_0# TEXT$20_0/m3_6480_0# 0
C1416 TEXT$21_0/m4_10080_0# TEXT$22_0/m2_10800_0# 0
C1417 TEXT$22_0/m2_9360_0# TEXT$1_0/m1_7200_0# 0
C1418 TEXT$21_0/m4_10800_0# TEXT$22_0/m2_10080_0# 0
C1419 TEXT$23_0/m1_14400_0# TEXT$6_0/m4_12000_0# -0
C1420 TEXT$3_0/m2_4800_0# TEXT$3_0/m2_6000_0# 0.20564f
C1421 PD VSS 2.34388f
C1422 VBIAS VSS 21.3749f
C1423 VIN VSS 21.5979f
C1424 VCM_OUT VSS 90.44077f
C1425 BCM_OUT VSS 83.53588f
C1426 CCM_OUT VSS 77.41045f
C1427 VIN_OUT VSS 75.9368f
C1428 TEXT$1_0/m1_12000_0# VSS 1.67051f
C1429 TEXT$1_0/m1_10800_0# VSS 1.57858f
C1430 TEXT$1_0/m1_9600_0# VSS 1.47068f
C1431 TEXT$1_0/m1_8400_0# VSS 1.61445f
C1432 TEXT$1_0/m1_7200_0# VSS 1.01495f
C1433 TEXT$1_0/m1_6000_0# VSS 1.47437f
C1434 TEXT$1_0/m1_4800_0# VSS 1.38135f
C1435 TEXT$1_0/m1_3600_0# VSS 1.50156f
C1436 TEXT$1_0/m1_2400_0# VSS 1.40096f
C1437 TEXT$1_0/m1_1200_0# VSS 1.47437f
C1438 TEXT$1_0/m1_0_0# VSS 1.55242f
C1439 M_0/a_410724_251737# VSS 2.90137f $ **FLOATING
C1440 M_0/a_410134_251737# VSS 7.50138f
C1441 M_0/a_409498_256643# VSS 9.69464f
C1442 M_0/a_409618_260539# VSS 8.70323f
C1443 M_0/a_404041_244568# VSS 14.12268f
C1444 M_0/a_403251_244568# VSS 6.25205f
C1445 M_0/a_402461_244568# VSS 9.17245f
C1446 a_498947_268180# VSS 0.20929p
C1447 M_0/a_404311_244568# VSS 0.16085f
C1448 M_0/a_403521_244568# VSS 0.03348f
C1449 M_0/a_402731_244568# VSS 0.03306f
C1450 M_0/a_401941_244568# VSS 0.03317f
C1451 M_0/a_401151_244568# VSS 2.63903f
C1452 m4_400150_261569# VSS 17.66492f
C1453 M_0/a_395162_259299# VSS 0.29295f $ **FLOATING
C1454 M_0/a_383940_262205# VSS 4.92556f $ **FLOATING
C1455 M_0/a_383620_262205# VSS 2.7563f $ **FLOATING
C1456 M_0/a_377450_262205# VSS 40.1477f $ **FLOATING
C1457 M_0/a_374398_259299# VSS 12.9247f $ **FLOATING
C1458 a_499016_248165# VSS 0.23231p
C1459 M_0/a_373878_259299# VSS 0.20081f $ **FLOATING
C1460 M_0/a_386992_259299# VSS 3.24772f $ **FLOATING
C1461 M_0/a_365708_259299# VSS 3.20723f $ **FLOATING
C1462 TEXT$3_0/m2_12000_0# VSS 1.10534f
C1463 TEXT$3_0/m2_10800_0# VSS 0.97985f
C1464 TEXT$3_0/m2_9600_0# VSS 0.92335f
C1465 TEXT$3_0/m2_8400_0# VSS 1.02903f
C1466 TEXT$3_0/m2_7200_0# VSS 0.67548f
C1467 TEXT$3_0/m2_6000_0# VSS 0.90425f
C1468 TEXT$3_0/m2_4800_0# VSS 0.84094f
C1469 TEXT$3_0/m2_3600_0# VSS 0.93809f
C1470 TEXT$3_0/m2_2400_0# VSS 0.86416f
C1471 TEXT$3_0/m2_1200_0# VSS 0.90425f
C1472 TEXT$3_0/m2_0_0# VSS 1.0227f
C1473 TEXT$21_0/m4_18000_0# VSS 0.3687f
C1474 TEXT$21_0/m4_17280_0# VSS 0.29292f
C1475 TEXT$21_0/m4_16560_0# VSS 0.25119f
C1476 TEXT$21_0/m4_15840_0# VSS 0.27618f
C1477 TEXT$21_0/m4_15120_0# VSS 0.26457f
C1478 TEXT$21_0/m4_14400_0# VSS 0.29187f
C1479 TEXT$21_0/m4_13680_0# VSS 0.25731f
C1480 TEXT$21_0/m4_12960_0# VSS 0.31454f
C1481 TEXT$21_0/m4_11700_0# VSS 0.17359f
C1482 TEXT$21_0/m4_10800_0# VSS 0.27936f
C1483 TEXT$21_0/m4_10080_0# VSS 0.29292f
C1484 TEXT$21_0/m4_9360_0# VSS 0.28243f
C1485 TEXT$21_0/m4_8640_0# VSS 0.28646f
C1486 TEXT$21_0/m4_7920_720# VSS 0.24565f
C1487 TEXT$21_0/m4_7200_0# VSS 0.27017f
C1488 TEXT$21_0/m4_6480_0# VSS 0.2796f
C1489 TEXT$21_0/m4_5760_0# VSS 0.31025f
C1490 TEXT$21_0/m4_4320_0# VSS 0.29779f
C1491 TEXT$21_0/m4_3780_0# VSS 0.15019f
C1492 TEXT$21_0/m4_2880_720# VSS 0.24684f
C1493 TEXT$21_0/m4_2160_0# VSS 0.27505f
C1494 TEXT$21_0/m4_1440_0# VSS 0.27946f
C1495 TEXT$21_0/m4_720_0# VSS 0.25389f
C1496 TEXT$21_0/m4_0_0# VSS 0.38208f
C1497 TEXT$23_0/m1_18000_0# VSS 0.74707f
C1498 TEXT$23_0/m1_17280_0# VSS 0.6816f
C1499 TEXT$23_0/m1_16560_0# VSS 0.60333f
C1500 TEXT$23_0/m1_15840_0# VSS 0.66424f
C1501 TEXT$23_0/m1_15120_0# VSS 0.63829f
C1502 TEXT$23_0/m1_14400_0# VSS 0.68975f
C1503 TEXT$23_0/m1_13680_0# VSS 0.61711f
C1504 TEXT$23_0/m1_12960_0# VSS 0.72574f
C1505 TEXT$23_0/m1_11700_0# VSS 0.43834f
C1506 TEXT$23_0/m1_10800_0# VSS 0.69166f
C1507 TEXT$23_0/m1_10080_0# VSS 0.6816f
C1508 TEXT$23_0/m1_9360_0# VSS 0.67042f
C1509 TEXT$23_0/m1_8640_0# VSS 0.7033f
C1510 TEXT$23_0/m1_7920_720# VSS 0.52865f
C1511 TEXT$23_0/m1_7200_0# VSS 0.62782f
C1512 TEXT$23_0/m1_6480_0# VSS 0.67466f
C1513 TEXT$23_0/m1_5760_0# VSS 0.72185f
C1514 TEXT$23_0/m1_4320_0# VSS 0.72911f
C1515 TEXT$23_0/m1_3780_0# VSS 0.40958f
C1516 TEXT$23_0/m1_2880_720# VSS 0.53649f
C1517 TEXT$23_0/m1_2160_0# VSS 0.68376f
C1518 TEXT$23_0/m1_1440_0# VSS 0.6748f
C1519 TEXT$23_0/m1_720_0# VSS 0.60668f
C1520 TEXT$23_0/m1_0_0# VSS 0.79623f
C1521 m3_419992_265695# VSS 0.1019p
C1522 EN VSS 6.16405f
C1523 TEXT$7_0/m2_10560_0# VSS 0.80673f
C1524 TEXT$7_0/m2_9600_0# VSS 0.73788f
C1525 TEXT$7_0/m2_7680_0# VSS 0.67937f
C1526 TEXT$7_0/m2_6720_0# VSS 0.66953f
C1527 TEXT$7_0/m2_5760_0# VSS 0.65242f
C1528 TEXT$7_0/m2_4800_960# VSS 0.50907f
C1529 TEXT$7_0/m2_3840_0# VSS 0.71466f
C1530 TEXT$7_0/m2_2880_0# VSS 0.62912f
C1531 TEXT$7_0/m2_2160_0# VSS 0.3654f
C1532 TEXT$7_0/m2_960_0# VSS 0.68878f
C1533 TEXT$7_0/m2_0_0# VSS 0.74409f
C1534 TEXT$9_0/m1_10560_0# VSS 1.21493f
C1535 TEXT$9_0/m1_9600_0# VSS 1.14824f
C1536 TEXT$9_0/m1_7680_0# VSS 1.05857f
C1537 TEXT$9_0/m1_6720_0# VSS 1.06655f
C1538 TEXT$9_0/m1_5760_0# VSS 1.04918f
C1539 TEXT$9_0/m1_4800_960# VSS 0.77249f
C1540 TEXT$9_0/m1_3840_0# VSS 1.14528f
C1541 TEXT$9_0/m1_2880_0# VSS 0.99494f
C1542 TEXT$9_0/m1_2160_0# VSS 0.60271f
C1543 TEXT$9_0/m1_960_0# VSS 1.09989f
C1544 TEXT$9_0/m1_0_0# VSS 1.09136f
C1545 TEXT$20_0/m3_18000_0# VSS 0.41838f
C1546 TEXT$20_0/m3_17280_0# VSS 0.34067f
C1547 TEXT$20_0/m3_16560_0# VSS 0.2941f
C1548 TEXT$20_0/m3_15840_0# VSS 0.32362f
C1549 TEXT$20_0/m3_15120_0# VSS 0.31056f
C1550 TEXT$20_0/m3_14400_0# VSS 0.34198f
C1551 TEXT$20_0/m3_13680_0# VSS 0.30197f
C1552 TEXT$20_0/m3_12960_0# VSS 0.36766f
C1553 TEXT$20_0/m3_11700_0# VSS 0.21174f
C1554 TEXT$20_0/m3_10800_0# VSS 0.33087f
C1555 TEXT$20_0/m3_10080_0# VSS 0.34067f
C1556 TEXT$20_0/m3_9360_0# VSS 0.32973f
C1557 TEXT$20_0/m3_8640_0# VSS 0.33785f
C1558 TEXT$20_0/m3_7920_720# VSS 0.2837f
C1559 TEXT$20_0/m3_7200_0# VSS 0.31599f
C1560 TEXT$20_0/m3_6480_0# VSS 0.32823f
C1561 TEXT$20_0/m3_5760_0# VSS 0.36291f
C1562 TEXT$20_0/m3_4320_0# VSS 0.35509f
C1563 TEXT$20_0/m3_3780_0# VSS 0.18429f
C1564 TEXT$20_0/m3_2880_720# VSS 0.28578f
C1565 TEXT$20_0/m3_2160_0# VSS 0.32657f
C1566 TEXT$20_0/m3_1440_0# VSS 0.3301f
C1567 TEXT$20_0/m3_720_0# VSS 0.29737f
C1568 TEXT$20_0/m3_0_0# VSS 0.43558f
C1569 TEXT$4_0/m3_12000_0# VSS 0.8798f
C1570 TEXT$4_0/m3_10800_0# VSS 0.74108f
C1571 TEXT$4_0/m3_9600_0# VSS 0.69952f
C1572 TEXT$4_0/m3_8400_0# VSS 0.78313f
C1573 TEXT$4_0/m3_7200_0# VSS 0.53411f
C1574 TEXT$4_0/m3_6000_0# VSS 0.68166f
C1575 TEXT$4_0/m3_4800_0# VSS 0.63268f
C1576 TEXT$4_0/m3_3600_0# VSS 0.71042f
C1577 TEXT$4_0/m3_2400_0# VSS 0.65181f
C1578 TEXT$4_0/m3_1200_0# VSS 0.68166f
C1579 TEXT$4_0/m3_0_0# VSS 0.81082f
C1580 TEXT$22_0/m2_18000_0# VSS 0.51369f
C1581 TEXT$22_0/m2_17280_0# VSS 0.43448f
C1582 TEXT$22_0/m2_16560_0# VSS 0.37855f
C1583 TEXT$22_0/m2_15840_0# VSS 0.41723f
C1584 TEXT$22_0/m2_15120_0# VSS 0.40122f
C1585 TEXT$22_0/m2_14400_0# VSS 0.43962f
C1586 TEXT$22_0/m2_13680_0# VSS 0.38971f
C1587 TEXT$22_0/m2_12960_0# VSS 0.46929f
C1588 TEXT$22_0/m2_11700_0# VSS 0.2813f
C1589 TEXT$22_0/m2_10800_0# VSS 0.4322f
C1590 TEXT$22_0/m2_10080_0# VSS 0.43448f
C1591 TEXT$22_0/m2_9360_0# VSS 0.42288f
C1592 TEXT$22_0/m2_8640_0# VSS 0.43926f
C1593 TEXT$22_0/m2_7920_720# VSS 0.35596f
C1594 TEXT$22_0/m2_7200_0# VSS 0.40444f
C1595 TEXT$22_0/m2_6480_0# VSS 0.42396f
C1596 TEXT$22_0/m2_5760_0# VSS 0.46439f
C1597 TEXT$22_0/m2_4320_0# VSS 0.4639f
C1598 TEXT$22_0/m2_3780_0# VSS 0.25019f
C1599 TEXT$22_0/m2_2880_720# VSS 0.36002f
C1600 TEXT$22_0/m2_2160_0# VSS 0.42722f
C1601 TEXT$22_0/m2_1440_0# VSS 0.42821f
C1602 TEXT$22_0/m2_720_0# VSS 0.38298f
C1603 TEXT$22_0/m2_0_0# VSS 0.53854f
C1604 TEXT$6_0/m4_12000_0# VSS 0.76245f
C1605 TEXT$6_0/m4_10800_0# VSS 0.61613f
C1606 TEXT$6_0/m4_9600_0# VSS 0.5809f
C1607 TEXT$6_0/m4_8400_0# VSS 0.65096f
C1608 TEXT$6_0/m4_7200_0# VSS 0.458f
C1609 TEXT$6_0/m4_6000_0# VSS 0.56715f
C1610 TEXT$6_0/m4_4800_0# VSS 0.5257f
C1611 TEXT$6_0/m4_3600_0# VSS 0.5906f
C1612 TEXT$6_0/m4_2400_0# VSS 0.54197f
C1613 TEXT$6_0/m4_1200_0# VSS 0.56715f
C1614 TEXT$6_0/m4_0_0# VSS 0.69997f
C1615 TEXT$24_0/m3_10560_0# VSS 0.66929f
C1616 TEXT$24_0/m3_9600_0# VSS 0.60631f
C1617 TEXT$24_0/m3_7680_0# VSS 0.53988f
C1618 TEXT$24_0/m3_6720_0# VSS 0.53604f
C1619 TEXT$24_0/m3_5760_0# VSS 0.50746f
C1620 TEXT$24_0/m3_4800_960# VSS 0.40695f
C1621 TEXT$24_0/m3_3840_0# VSS 0.55397f
C1622 TEXT$24_0/m3_2880_0# VSS 0.48843f
C1623 TEXT$24_0/m3_2160_0# VSS 0.28113f
C1624 TEXT$24_0/m3_960_0# VSS 0.53366f
C1625 TEXT$24_0/m3_0_0# VSS 0.62072f
C1626 TEXT$8_0/m4_10560_0# VSS 0.58619f
C1627 TEXT$8_0/m4_9600_0# VSS 0.52311f
C1628 TEXT$8_0/m4_7680_0# VSS 0.46028f
C1629 TEXT$8_0/m4_6720_0# VSS 0.45506f
C1630 TEXT$8_0/m4_5760_0# VSS 0.42745f
C1631 TEXT$8_0/m4_4800_960# VSS 0.35093f
C1632 TEXT$8_0/m4_3840_0# VSS 0.46517f
C1633 TEXT$8_0/m4_2880_0# VSS 0.41267f
C1634 TEXT$8_0/m4_2160_0# VSS 0.23197f
C1635 TEXT$8_0/m4_960_0# VSS 0.44746f
C1636 TEXT$8_0/m4_0_0# VSS 0.54263f
C1637 VDD VSS 2.42752p
C1638 PU VSS 5.85351f
C1639 sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tiel$3_0/a_124_157# VSS 0.3723f
C1640 sc_tieh_tiel$1_0/gf180mcu_fd_sc_mcu9t5v0__tieh$2_0/a_125_157# VSS 0.37323f
.ends

