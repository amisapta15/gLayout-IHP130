** sch_path: /foss/pdks/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/tran_logic_nand.sch
**.subckt tran_logic_nand
VinA A GND dc 0 ac 0 pulse(0, 1.2, 2n, 100p, 100p, 4n, 6n )
Vdd net1 GND 1.2
VinB B GND dc 0 ac 0 pulse(0, 1.2, 0, 100p, 100p, 2n, 4n )
XM1 net2 A GND GND sg13_lv_nmos w=1.0u l=0.45u ng=1 m=1
XM3 out B net2 GND sg13_lv_nmos w=1.0u l=0.45u ng=1 m=1
XM2 out A net1 net1 sg13_lv_pmos w=1.0u l=0.45u ng=1 m=1
XM4 out B net1 net1 sg13_lv_pmos w=1.0u l=0.45u ng=1 m=1
**** begin user architecture code

.lib cornerMOSlv.lib mos_ff



.param temp=127
.control
save all
tran 50p 20n
meas tran tdelay TRIG v(b) VAl=0.9 FALl=1 TARG v(out) VAl=0.9 RISE=1
write tran_logic_nand.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
