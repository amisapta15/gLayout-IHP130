** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/trimmer.sch
**.subckt trimmer
XMP1 net1 net1 VDD VDD sg13_lv_pmos w=0.28u l=8.0u ng=1 m=1
XMP2 net2 net2 net1 VDD sg13_lv_pmos w=0.28u l=8.0u ng=1 m=1
XMN2 net4 net2 GND GND sg13_lv_nmos w=0.28u l=8.0u ng=1 m=1
XMN1 net2 net2 GND GND sg13_lv_nmos w=0.28u l=8.0u ng=1 m=1
XMP3 net3 net5 VDD VDD sg13_lv_pmos w=2.0u l=2.0u ng=2 m=1
XMP4 net4 VDD net3 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP5 net6 net5 VDD VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=2
XMP6 net8 VDD net6 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP7 net7 net5 VDD VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=2
XMP8 vbp VDD net7 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP9 net8 net4 VDD VDD sg13_lv_pmos w=0.28u l=8.0u ng=1 m=1
XMN3 net8 net8 GND GND sg13_lv_nmos w=2.0u l=2.0u ng=1 m=1
XMN4 vbp_casc net8 net9 GND sg13_lv_nmos w=2.0u l=2.0u ng=1 m=4
XR1 vbp_casc vbp sub! rppd w=0.5e-6 l=389e-6 m=1 b=0
XR2 GND net9 sub! rhigh w=0.5e-6 l=152.5e-6 m=1 b=0
vbp net5 vbp 0
.save i(vbp)
vbp_casc VDD vbp_casc 0
.save i(vbp_casc)
Vdd VDD GND 1.8
R3 net13 net14 300 m=1
XMP10 net10 vbp VDD VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=2
XMP11 net13 vbp_casc net10 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP12 net11 vbp net15 VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=4
XMP13 net13 vbp_casc net11 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=4
XMP14 net12 vbp net16 VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=8
XMP15 net13 vbp_casc net12 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=8
vload net14 GND 0
.save i(vload)
**** begin user architecture code


* --- parameters ---
.param Rload = 300
.control
  set noaskquit
  step param Rload list 50 100 150 200 300
  op
  plot Rload vs i(vload)
.endc



 .lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ_stat

**** end user architecture code
**.ends
.GLOBAL GND
.end
