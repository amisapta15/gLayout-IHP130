** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/DPI_try_1.sch
**.subckt DPI_try_1
Vgs G GND -0.75
Vds D GND -1.5
Vd D net1 0
.save i(vd)
XM3 net1 G GND GND sg13_lv_pmos w=1.0u l=0.45u ng=1 m=1
**** begin user architecture code


.options savecurrrents
.include DPI_try_1.save
.param temp=27
.control
save all
op
write DPI_try_1.raw
set appendwrite
*dc Vds 0 1.2 0.01 Vgs 0.3 1.0 0.1
*dc Vgs 0 0.5 0.05
dc vds 0 -1.2 -0.01 Vgs -0.35 -1.1 -0.05
write DPI_try_1.raw
.endc


 .lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
