| units: 0.5 tech: gf180mcuD format: MIT
x a_n1900_n6686# VDD a_n1900_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1779 y=-1337 pfet_03v3
x a_n28653_8045# a_n25601_10951# a_n28653_8045# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-23120 y=10951 nfet_03v3
x VIN a_470_n6686# a_990_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=590 y=-6685 pfet_03v3
x EN VDD a_n1900_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=195 y=4114 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=6595 y=-1654 nfet_03v3
x VSS VSS VSS VSS d=185600,3432 l=200 w=1600 x=-18702 y=10951 nfet_03v3
x a_990_n6686# VSS a_6447_5389# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7157 y=7527 nfet_03v3
x a_n37343_8045# VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-36432 y=10951 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-28244 y=8045 pfet_03v3
x a_7083_483# VSS a_7083_483# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7203 y=-1654 nfet_03v3
x a_990_n6686# VSS a_6447_5389# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=8337 y=7527 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=2188 y=-6685 pfet_03v3
x VAUX a_n37343_8045# VAUX VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-33272 y=8045 pfet_03v3
x a_n16059_8045# VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-13568 y=10951 pfet_03v3
x a_n25601_10951# VSS a_n25601_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-23120 y=8445 nfet_03v3
x a_n19111_10951# a_n16059_8045# a_n19111_10951# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-8828 y=8045 pfet_03v3
x a_n25601_10951# VSS a_n25601_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-24300 y=8445 nfet_03v3
x a_n28653_8045# a_n25601_10951# a_n28653_8045# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-21350 y=10951 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-28244 y=10951 pfet_03v3
x VAUX a_n37343_8045# VAUX VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-34852 y=8045 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=6595 y=483 nfet_03v3
x VSS VSS VSS VSS d=185600,3432 l=200 w=1600 x=-26088 y=10951 nfet_03v3
x VIN a_n1110_n6686# a_n590_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-989 y=-6685 pfet_03v3
x a_n19111_10951# a_n16059_8045# a_n19111_10951# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-13568 y=8045 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2587 y=-6685 pfet_03v3
x EN VDD a_n1900_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-594 y=4114 pfet_03v3
x EN VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-15938 y=14649 pfet_03v3
x a_n28653_8045# a_n25601_10951# a_n28653_8045# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-25480 y=10951 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=6595 y=-8696 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2192 y=4114 pfet_03v3
x a_n25601_10951# VSS a_n25601_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-24890 y=8445 nfet_03v3
x VAUX a_n37343_8045# VAUX VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-37222 y=8045 pfet_03v3
x VSS VSS VSS VSS d=185600,3432 l=200 w=1600 x=-26088 y=8445 nfet_03v3
x a_n37343_8045# VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-34852 y=10951 pfet_03v3
x a_n19111_10951# a_n7889_8045# a_n7369_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-7768 y=8045 pfet_03v3
x EN VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-37222 y=14649 pfet_03v3
x a_n590_n6686# VSS a_n590_n6686# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7203 y=-8696 nfet_03v3
x a_n28653_8045# a_n25601_10951# a_n28653_8045# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-24300 y=10951 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5959 y=5389 nfet_03v3
x a_n16059_8045# VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-11988 y=10951 pfet_03v3
x VSS VSS VSS VSS d=185600,3432 l=200 w=1600 x=-18702 y=8445 nfet_03v3
x a_n1900_n6686# VDD a_470_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=590 y=-1337 pfet_03v3
x a_n37343_8045# VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-33272 y=10951 pfet_03v3
x VIN a_1260_n6686# VOUT_VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=1380 y=-6685 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-15130 y=14649 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8945 y=5389 nfet_03v3
x EN VDD a_n1900_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=985 y=4114 pfet_03v3
x a_n7369_8045# a_6447_5389# VOUT_RCCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6567 y=5389 nfet_03v3
x a_n25601_10951# VSS a_n19431_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-19310 y=8445 nfet_03v3
x VAUX a_n37343_8045# VAUX VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-32482 y=8045 pfet_03v3
x VAUX a_n37343_8045# VAUX VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-30112 y=8045 pfet_03v3
x a_n7369_8045# a_6447_5389# VOUT_RCCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7747 y=5389 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=2188 y=-1337 pfet_03v3
x a_n25601_10951# VSS a_n25601_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-25480 y=8445 nfet_03v3
x a_7083_483# VSS a_7673_483# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7793 y=-1654 nfet_03v3
x a_n16059_8045# VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-15938 y=10951 pfet_03v3
x a_n28653_8045# a_n25601_10951# a_n28653_8045# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-22530 y=10951 nfet_03v3
x a_n19111_10951# a_n16059_8045# a_n19111_10951# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-11198 y=8045 pfet_03v3
x a_n37343_8045# VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-37222 y=10951 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8401 y=-1654 nfet_03v3
x a_n37343_8045# VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-30902 y=10951 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5959 y=9665 nfet_03v3
x a_n19111_10951# a_n16059_8045# a_n19111_10951# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-12778 y=8045 pfet_03v3
x a_n1900_n6686# VDD a_n1110_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-989 y=-1337 pfet_03v3
x a_n19111_10951# a_n16059_8045# a_n19111_10951# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-10408 y=8045 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2587 y=-1337 pfet_03v3
x a_n16059_8045# VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-8828 y=10951 pfet_03v3
x a_n16059_8045# VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-14358 y=10951 pfet_03v3
x a_n37343_8045# VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-31692 y=10951 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8945 y=9665 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-16746 y=8045 pfet_03v3
x VAUX a_n37343_8045# VAUX VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-36432 y=8045 pfet_03v3
x a_n28653_8045# a_n25601_10951# a_n28653_8045# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-20760 y=10951 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8401 y=483 nfet_03v3
x a_6447_5389# VSS a_n7369_8045# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7157 y=5389 nfet_03v3
x a_n19111_10951# a_n16059_8045# a_n19111_10951# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-15148 y=8045 pfet_03v3
x a_6567_9285# VSS a_n7369_8045# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6567 y=9665 nfet_03v3
x a_6447_5389# VSS a_n7369_8045# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=8337 y=5389 nfet_03v3
x a_6567_9285# VSS a_n7369_8045# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7747 y=9665 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1793 y=4114 pfet_03v3
x a_n590_n6686# VSS VOUT_VCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7793 y=-8696 nfet_03v3
x EN VDD a_n1900_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1384 y=4114 pfet_03v3
x a_n28653_8045# a_n25601_10951# a_n28653_8045# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-24890 y=10951 nfet_03v3
x a_n1900_n6686# VDD a_1260_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=1380 y=-1337 pfet_03v3
x a_n16059_8045# VDD a_n7889_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-7768 y=10951 pfet_03v3
x a_n37343_8045# VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-35642 y=10951 pfet_03v3
x VAUX a_n29173_8045# a_n28653_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-29052 y=8045 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8401 y=-8696 nfet_03v3
x a_n37343_8045# VDD a_n29173_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-29052 y=10951 pfet_03v3
x VIN a_n320_n6686# a_200_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-199 y=-6685 pfet_03v3
x VIN a_n1900_n6686# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1779 y=-6685 pfet_03v3
x a_n16059_8045# VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-12778 y=10951 pfet_03v3
x a_n28653_8045# a_n25601_10951# a_n28653_8045# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-23710 y=10951 nfet_03v3
x VAUX a_n37343_8045# VAUX VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-31692 y=8045 pfet_03v3
x a_n16059_8045# VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-10408 y=10951 pfet_03v3
x a_n25601_10951# VSS a_n25601_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-20760 y=8445 nfet_03v3
x a_n28653_8045# a_n19431_10951# a_n19111_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-19310 y=10951 nfet_03v3
x a_n37343_8045# VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-34062 y=10951 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-16746 y=14649 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-36414 y=14649 pfet_03v3
x a_n25601_10951# VSS a_n25601_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-21940 y=8445 nfet_03v3
x a_200_n6686# a_7083_483# a_200_n6686# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7203 y=483 nfet_03v3
x a_n7369_8045# a_6567_9285# a_990_n6686# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7157 y=9665 nfet_03v3
x VAUX a_n37343_8045# VAUX VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-30902 y=8045 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5959 y=7527 nfet_03v3
x a_n7369_8045# a_6567_9285# a_990_n6686# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=8337 y=9665 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-38030 y=14649 pfet_03v3
x a_n16059_8045# VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-11198 y=10951 pfet_03v3
x a_n19111_10951# a_n16059_8045# a_n19111_10951# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-11988 y=8045 pfet_03v3
x VAUX a_n37343_8045# VAUX VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-34062 y=8045 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8945 y=7527 nfet_03v3
x a_n19111_10951# a_n16059_8045# a_n19111_10951# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-9618 y=8045 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-38030 y=8045 pfet_03v3
x a_n28653_8045# a_n25601_10951# a_n28653_8045# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-21940 y=10951 nfet_03v3
x VAUX a_n37343_8045# VAUX VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-35642 y=8045 pfet_03v3
x a_990_n6686# VSS a_6567_9285# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6567 y=7527 nfet_03v3
x a_n28653_8045# a_n25601_10951# a_n28653_8045# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-20170 y=10951 nfet_03v3
x a_n19111_10951# a_n16059_8045# a_n19111_10951# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-14358 y=8045 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-6960 y=10951 pfet_03v3
x a_990_n6686# VSS a_6567_9285# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7747 y=7527 nfet_03v3
x a_n25601_10951# VSS a_n25601_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-20170 y=8445 nfet_03v3
x a_n16059_8045# VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-9618 y=10951 pfet_03v3
x a_n16059_8045# VDD a_n16059_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-15148 y=10951 pfet_03v3
x a_n25601_10951# VSS a_n25601_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-21350 y=8445 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-6960 y=8045 pfet_03v3
x a_n19111_10951# a_n16059_8045# a_n19111_10951# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-15938 y=8045 pfet_03v3
x a_n37343_8045# VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-32482 y=10951 pfet_03v3
x a_n25601_10951# VSS a_n25601_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-22530 y=8445 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-16746 y=10951 pfet_03v3
x a_n37343_8045# VDD a_n37343_8045# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-30112 y=10951 pfet_03v3
x a_n25601_10951# VSS a_n25601_10951# VSS s=192000,3440 d=192000,3440 l=200 w=1600 x=-23710 y=8445 nfet_03v3
x a_200_n6686# a_7673_483# VOUT_SBCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7793 y=483 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-38030 y=10951 pfet_03v3
x a_n1900_n6686# VDD a_n320_n6686# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-199 y=-1337 pfet_03v3
C a_n29173_8045# VAUX 1.0
C a_1260_n6686# a_470_n6686# 0.8
C EN a_470_n6686# 0.0
C a_7673_483# a_7083_483# 0.4
C a_n1110_n6686# VIN 2.9
C a_990_n6686# VIN 0.6
C VOUT_VIN a_470_n6686# 0.1
C a_n7889_8045# VDD 3.1
C a_n590_n6686# VIN 0.6
C a_1260_n6686# a_200_n6686# 0.1
C a_n19111_10951# a_n16059_8045# 29.5
C a_n28653_8045# EN 0.0
C VDD a_470_n6686# 7.5
C a_200_n6686# VOUT_VIN 0.1
C VOUT_RCCM a_6567_9285# 0.0
C a_n25601_10951# a_n19431_10951# 0.5
C a_n37343_8045# a_n28653_8045# 0.1
C VDD a_200_n6686# 1.1
C a_6567_9285# a_6447_5389# 0.4
C a_1260_n6686# a_n1110_n6686# 0.3
C a_n28653_8045# VDD 1.8
C EN a_n19111_10951# 0.0
C a_990_n6686# a_1260_n6686# 2.3
C a_1260_n6686# a_n590_n6686# 0.1
C EN a_n1110_n6686# 0.0
C EN a_n29173_8045# 0.0
C a_n1110_n6686# VOUT_VIN 0.1
C a_990_n6686# VOUT_VIN 2.5
C a_n590_n6686# VOUT_VIN 0.1
C a_n37343_8045# a_n29173_8045# 1.0
C a_n19111_10951# VDD 15.5
C VDD a_n1110_n6686# 7.4
C a_n1900_n6686# a_n320_n6686# 1.5
C a_990_n6686# VDD 1.7
C a_7673_483# VOUT_SBCM 1.2
C VDD a_n29173_8045# 3.1
C a_990_n6686# a_6567_9285# 3.0
C a_200_n6686# a_470_n6686# 2.3
C a_n590_n6686# VDD 1.2
C VOUT_SBCM a_7083_483# 0.1
C VOUT_RCCM a_6447_5389# 2.2
C a_n19111_10951# a_n7889_8045# 1.0
C a_n16059_8045# a_n7369_8045# 0.1
C VIN a_n320_n6686# 0.6
C a_n1110_n6686# a_470_n6686# 0.3
C a_990_n6686# a_470_n6686# 2.4
C a_n590_n6686# a_470_n6686# 0.1
C a_990_n6686# VOUT_RCCM 0.0
C a_n1900_n6686# VIN 3.4
C a_200_n6686# a_n1110_n6686# 0.2
C EN a_n7369_8045# 0.0
C a_n28653_8045# a_n19111_10951# 0.3
C VAUX VIN 0.0
C a_990_n6686# a_200_n6686# 0.3
C a_990_n6686# a_6447_5389# 0.9
C a_n590_n6686# a_200_n6686# 0.6
C a_n28653_8045# a_n29173_8045# 0.9
C a_n7369_8045# VOUT_VIN 0.2
C a_1260_n6686# a_n320_n6686# 0.3
C a_n590_n6686# VOUT_VCM 0.2
C EN a_n320_n6686# 0.0
C VOUT_SBCM VIN 0.1
C a_n320_n6686# VOUT_VIN 0.1
C VDD a_n7369_8045# 1.6
C a_n7369_8045# a_6567_9285# 3.6
C a_n1900_n6686# a_1260_n6686# 2.4
C a_990_n6686# a_n1110_n6686# 0.2
C a_n590_n6686# a_n1110_n6686# 2.4
C EN a_n1900_n6686# 2.2
C a_990_n6686# a_n590_n6686# 0.1
C VDD a_n320_n6686# 7.4
C a_n1900_n6686# VOUT_VIN 1.0
C a_n7889_8045# a_n7369_8045# 0.9
C EN VAUX 0.0
C a_n25601_10951# a_n28653_8045# 36.6
C a_1260_n6686# VIN 0.6
C a_n1900_n6686# VDD 44.9
C EN VIN 0.1
C a_n37343_8045# VAUX 29.5
C VOUT_RCCM a_n7369_8045# 0.6
C a_7673_483# a_200_n6686# 1.5
C VIN VOUT_VIN 0.6
C VDD VAUX 16.3
C a_200_n6686# a_7083_483# 1.9
C a_n320_n6686# a_470_n6686# 0.8
C EN a_n16059_8045# 0.8
C a_n7369_8045# a_6447_5389# 3.3
C VDD VIN 14.6
C a_200_n6686# a_n320_n6686# 2.4
C a_n1900_n6686# a_470_n6686# 1.5
C a_n16059_8045# VDD 48.8
C EN a_1260_n6686# 0.3
C a_n19111_10951# a_n7369_8045# 0.5
C a_1260_n6686# VOUT_VIN 2.4
C a_990_n6686# a_n7369_8045# 1.5
C a_n1900_n6686# a_200_n6686# 0.1
C VIN a_470_n6686# 0.6
C a_n7889_8045# a_n16059_8045# 1.0
C a_n37343_8045# EN 0.7
C a_n1110_n6686# a_n320_n6686# 0.8
C a_1260_n6686# VDD 6.4
C VOUT_RCCM VIN 0.1
C a_n28653_8045# a_n19431_10951# 0.9
C a_990_n6686# a_n320_n6686# 0.2
C a_n28653_8045# VAUX 0.5
C a_n590_n6686# a_n320_n6686# 2.3
C EN VDD 19.3
C VDD VOUT_VIN 2.9
C a_6567_9285# VOUT_VIN 0.0
C a_200_n6686# VIN 0.6
C VOUT_SBCM a_200_n6686# 0.2
C a_n1900_n6686# a_n1110_n6686# 1.8
C VOUT_VCM VIN 0.1
C a_n37343_8045# VDD 48.9
C a_990_n6686# a_n1900_n6686# 0.6
C a_n1900_n6686# a_n590_n6686# 0.1
C EN a_n7889_8045# 0.0
C a_n19111_10951# a_n19431_10951# 1.1
C VOUT_VCM0 6.1
R VOUT_VCM 55
C VOUT_SBCM0 4.7
R VOUT_SBCM 55
C VOUT_RCCM0 6.0
R VOUT_RCCM 114
C VOUT_VIN0 10.5
R VOUT_VIN 154
C VIN0 33.1
R VIN 573
C VAUX0 25.4
R VAUX 2060
C EN0 24.1
R EN 462
C VDD0 950.0
R VDD 38605
R VSS 12140
C a_7673_483#0 2.9
R a_7673_483# 107
C a_7083_483#0 6.4
R a_7083_483# 219
C a_6447_5389#0 8.5
R a_6447_5389# 340
C a_6567_9285#0 7.7
R a_6567_9285# 335
C a_990_n6686#0 11.5
R a_990_n6686# 489
C a_200_n6686#0 5.1
R a_200_n6686# 293
C a_n590_n6686#0 8.0
R a_n590_n6686# 292
C a_1260_n6686#0 0.2
R a_1260_n6686# 272
C a_470_n6686#0 0.0
R a_470_n6686# 272
C a_n320_n6686#0 0.0
R a_n320_n6686# 272
C a_n1110_n6686#0 0.0
R a_n1110_n6686# 272
C a_n1900_n6686#0 2.6
R a_n1900_n6686# 1220
C a_n7369_8045#0 18.2
R a_n7369_8045# 603
C a_n7889_8045#0 0.3
R a_n7889_8045# 260
C a_n19111_10951#0 4.9
R a_n19111_10951# 2090
C a_n19431_10951#0 2.8
R a_n19431_10951# 191
C a_n25601_10951#0 40.1
R a_n25601_10951# 2962
C a_n28653_8045#0 12.9
R a_n28653_8045# 2054
C a_n29173_8045#0 0.2
R a_n29173_8045# 260
C a_n16059_8045#0 3.2
R a_n16059_8045# 3505
C a_n37343_8045#0 3.2
R a_n37343_8045# 3505
