** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/trimmer.sch
**.subckt trimmer
XMP1 net1 net1 net12 VDD sg13_lv_pmos w=0.28u l=8.0u ng=1 m=1
XMP2 vstart vstart net1 VDD sg13_lv_pmos w=0.28u l=8.0u ng=1 m=1
XMN2 net3 vstart GND GND sg13_lv_nmos w=0.28u l=8.0u ng=1 m=1
XMN1 vstart vstart GND GND sg13_lv_nmos w=0.28u l=8.0u ng=1 m=1
XMP3 net2 vbp net11 VDD sg13_lv_pmos w=2.0u l=2.0u ng=2 m=1
XMP4 net3 vbp_casc net2 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP5 net4 vbp net10 VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=2
XMP6 net6 vbp_casc net4 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP7 net5 vbp net9 VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=2
XMP8 vbp vbp_casc net5 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP9 net6 net3 enN VDD sg13_lv_pmos w=0.28u l=8.0u ng=1 m=1
XMN3 net6 net6 GND GND sg13_lv_nmos w=2.0u l=2.0u ng=1 m=1
XMN4 vbp_casc net6 net7 GND sg13_lv_nmos w=2.0u l=2.0u ng=1 m=4
XR1 vbp_casc vbp rppd w=0.5e-6 l=389e-6 m=1 b=0
XR2 GND net7 rhigh w=0.5e-6 l=152.5e-6 m=1 b=0
R3 ibias GND 300 m=1
XMP10 net8 vbp VDD VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=2
XMP11 ibias vbp_casc net8 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP16 vbp_casc enMon VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=1
XMP17 net9 enN VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=1
XMP18 net10 enN VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=1
XMP19 net12 enN VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=1
XMP20 net11 enN VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=1
XMN5 vstart enN GND GND sg13_lv_nmos w=2u l=0.28u ng=1 m=1
XMN6 net6 enN GND GND sg13_lv_nmos w=2u l=0.28u ng=1 m=1
V1 VDD GND 1.65
Ven en GND 1.65
xinv1 VDD en enN GND inv
xinv2 VDD enN enMon GND inv
XMP12 net13 vbp VDD VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=4
XMP13 ibias vbp_casc net13 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP14 net14 vbp VDD VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=8
XMP15 ibias vbp_casc net14 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
**** begin user architecture code


.include trimmer.save
.option savecurrent
.param temp=127
.control
op
save all
tran 500p 65u
plot en enN enMon
plot vstart
plot vbp vbp_casc
plot v(ibias)/300
.endc





.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ


**** end user architecture code
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/inv.sym
** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/inv.sch
.subckt inv VDD in out VSS
*.iopin VDD
*.ipin in
*.iopin VSS
*.opin out
XM1 out in VSS VSS sg13_lv_nmos w=2.0u l=0.28u ng=1 m=1
XM2 out in VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=1
.ends

.GLOBAL GND
.end
