* NGSPICE file created from M.ext - technology: gf180mcuD

.subckt M VIN VSS VDD VOUT_VIN VOUT_RCCM VOUT_SBCM VOUT_VCM VAUX EN
X0 a_n1900_n6686# a_n1900_n6686# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X1 a_n28653_8045# a_n28653_8045# a_n25601_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X2 a_990_n6686# VIN a_470_n6686# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X3 a_n1900_n6686# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X4 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0.1744n ps=0.65672m w=4u l=1u
X5 VSS VSS VSS VSS nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X6 a_6447_5389# a_990_n6686# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X7 a_n37343_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X8 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0.4068n ps=1.46136m w=10u l=2u
X9 a_7083_483# a_7083_483# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X10 a_6447_5389# a_990_n6686# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X11 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X12 VAUX VAUX a_n37343_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X13 a_n16059_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X14 a_n25601_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X15 a_n19111_10951# a_n19111_10951# a_n16059_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X16 a_n25601_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X17 a_n28653_8045# a_n28653_8045# a_n25601_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X18 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X19 VAUX VAUX a_n37343_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X20 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X21 VSS VSS VSS VSS nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X22 a_n590_n6686# VIN a_n1110_n6686# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X23 a_n19111_10951# a_n19111_10951# a_n16059_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X24 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X25 a_n1900_n6686# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X26 a_n16059_8045# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X27 a_n28653_8045# a_n28653_8045# a_n25601_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X28 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X29 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X30 a_n25601_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X31 VAUX VAUX a_n37343_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X32 VSS VSS VSS VSS nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X33 a_n37343_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X34 a_n7369_8045# a_n19111_10951# a_n7889_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X35 a_n37343_8045# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X36 a_n590_n6686# a_n590_n6686# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X37 a_n28653_8045# a_n28653_8045# a_n25601_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X38 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X39 a_n16059_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X40 VSS VSS VSS VSS nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X41 a_470_n6686# a_n1900_n6686# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X42 a_n37343_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X43 VOUT_VIN VIN a_1260_n6686# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X44 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X45 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X46 a_n1900_n6686# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X47 VOUT_RCCM a_n7369_8045# a_6447_5389# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X48 a_n19431_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X49 VAUX VAUX a_n37343_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X50 VAUX VAUX a_n37343_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X51 VOUT_RCCM a_n7369_8045# a_6447_5389# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X52 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X53 a_n25601_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X54 a_7673_483# a_7083_483# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X55 a_n16059_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X56 a_n28653_8045# a_n28653_8045# a_n25601_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X57 a_n19111_10951# a_n19111_10951# a_n16059_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X58 a_n37343_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X59 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X60 a_n37343_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X61 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X62 a_n19111_10951# a_n19111_10951# a_n16059_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X63 a_n1110_n6686# a_n1900_n6686# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X64 a_n19111_10951# a_n19111_10951# a_n16059_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X65 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X66 a_n16059_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X67 a_n16059_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X68 a_n37343_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X69 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X70 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X71 VAUX VAUX a_n37343_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X72 a_n28653_8045# a_n28653_8045# a_n25601_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X73 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X74 a_n7369_8045# a_6447_5389# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X75 a_n19111_10951# a_n19111_10951# a_n16059_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X76 a_n7369_8045# a_6567_9285# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X77 a_n7369_8045# a_6447_5389# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X78 a_n7369_8045# a_6567_9285# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X79 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X80 VOUT_VCM a_n590_n6686# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X81 a_n1900_n6686# EN VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X82 a_n28653_8045# a_n28653_8045# a_n25601_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X83 a_1260_n6686# a_n1900_n6686# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X84 a_n7889_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X85 a_n37343_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X86 a_n28653_8045# VAUX a_n29173_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X87 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X88 a_n29173_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X89 a_200_n6686# VIN a_n320_n6686# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X90 VIN VIN a_n1900_n6686# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X91 a_n16059_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X92 a_n28653_8045# a_n28653_8045# a_n25601_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X93 VAUX VAUX a_n37343_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X94 a_n16059_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X95 a_n25601_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X96 a_n19111_10951# a_n28653_8045# a_n19431_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X97 a_n37343_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X98 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X99 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X100 a_n25601_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X101 a_200_n6686# a_200_n6686# a_7083_483# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X102 a_990_n6686# a_n7369_8045# a_6567_9285# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X103 VAUX VAUX a_n37343_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X104 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X105 a_990_n6686# a_n7369_8045# a_6567_9285# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X106 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X107 a_n16059_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X108 a_n19111_10951# a_n19111_10951# a_n16059_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X109 VAUX VAUX a_n37343_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X110 VSS VSS VSS VSS nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X111 a_n19111_10951# a_n19111_10951# a_n16059_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X112 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X113 a_n28653_8045# a_n28653_8045# a_n25601_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X114 VAUX VAUX a_n37343_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X115 a_6567_9285# a_990_n6686# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X116 a_n28653_8045# a_n28653_8045# a_n25601_10951# VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X117 a_n19111_10951# a_n19111_10951# a_n16059_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X118 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X119 a_6567_9285# a_990_n6686# VSS VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X120 a_n25601_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X121 a_n16059_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X122 a_n16059_8045# a_n16059_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X123 a_n25601_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X124 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X125 a_n19111_10951# a_n19111_10951# a_n16059_8045# VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X126 a_n37343_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X127 a_n25601_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X128 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X129 a_n37343_8045# a_n37343_8045# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X130 a_n25601_10951# a_n25601_10951# VSS VSS nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X131 VOUT_SBCM a_200_n6686# a_7673_483# VSS nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X132 VDD VDD VDD VDD pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X133 a_n320_n6686# a_n1900_n6686# VDD VDD pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
.ends

