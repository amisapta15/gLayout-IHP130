** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/block_1_input.sch
**.subckt block_1_input
XM6 net1 net1 VDD VDD sg13_lv_pmos w=1.0u l=0.45u ng=1 m=1
XM7 net2 net1 VDD VDD sg13_lv_pmos w=1.0u l=0.45u ng=1 m=1
Icop net2 net4 0
.save i(icop)
Vdd VDD GND 1.2
I0 VDD net3 pulse(0 10n 0 1n 1n 10n 20n)
Iin net3 net1 0
.save i(iin)
VIn net4 GND 0
**** begin user architecture code



.options savecurrents
.include block_1_input.save

.param temp=27
.control
save all

op

write block_1_input.raw
set appendwrite

tran 1p 100n

plot i(VIn)

write block_1_input.raw
.endc


 .lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
