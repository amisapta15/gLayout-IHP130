* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu9t5v0__tieh$2 VDD VSS Z VNW VPW
X0 Z a_125_157# VDD VNW pfet_05v0 ad=0.396p pd=2.68u as=0.396p ps=2.68u w=0.9u l=0.5u
X1 a_125_157# a_125_157# VSS VPW nfet_05v0 ad=0.2904p pd=2.2u as=0.2904p ps=2.2u w=0.66u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__tiel$3 VDD VSS ZN VNW VPW
X0 ZN a_124_157# VSS VPW nfet_05v0 ad=0.2904p pd=2.2u as=0.2904p ps=2.2u w=0.66u l=0.6u
X1 a_124_157# a_124_157# VDD VNW pfet_05v0 ad=0.396p pd=2.68u as=0.396p ps=2.68u w=0.9u l=0.5u
.ends

.subckt sc_tieh_tiel$1 tieH tieL VDD VSS
Xgf180mcu_fd_sc_mcu9t5v0__tieh$2_0 VDD VSS tieH VDD VSS gf180mcu_fd_sc_mcu9t5v0__tieh$2
Xgf180mcu_fd_sc_mcu9t5v0__tiel$3_0 VDD VSS tieL VDD VSS gf180mcu_fd_sc_mcu9t5v0__tiel$3
.ends

.subckt ppolyf_u_9H3LNU$2 a_n224793_504053# w_n225009_503837# a_n224793_506155#
X0 a_n224793_506155# a_n224793_504053# w_n225009_503837# ppolyf_u r_width=40u r_length=10u
.ends

.subckt diode_nd2ps_06v0_MV3SZ3$2 a_505271_219793# a_503039_219793# a_507503_219793#
+ a_500807_219793# a_500655_219641#
D0 a_500655_219641# a_505271_219793# diode_nd2ps_06v0 pj=40u area=99.99999p
D1 a_500655_219641# a_500807_219793# diode_nd2ps_06v0 pj=40u area=99.99999p
D2 a_500655_219641# a_503039_219793# diode_nd2ps_06v0 pj=40u area=99.99999p
D3 a_500655_219641# a_507503_219793# diode_nd2ps_06v0 pj=40u area=99.99999p
.ends

.subckt diode_pd2nw_06v0_5DG9HC$2 a_507479_219793# a_500831_219793# w_500655_219617#
+ a_503047_219793# a_505263_219793#
D0 a_500831_219793# w_500655_219617# diode_pd2nw_06v0 pj=40u area=99.99999p
D1 a_507479_219793# w_500655_219617# diode_pd2nw_06v0 pj=40u area=99.99999p
D2 a_503047_219793# w_500655_219617# diode_pd2nw_06v0 pj=40u area=99.99999p
D3 a_505263_219793# w_500655_219617# diode_pd2nw_06v0 pj=40u area=99.99999p
.ends

.subckt io_secondary_5p0$1 m1_499212_228525# m1_497955_232243# m1_512035_219553# VSUBS
Xppolyf_u_9H3LNU_0 m1_499212_228525# m1_497955_232243# m1_512035_219553# ppolyf_u_9H3LNU$2
Xdiode_nd2ps_06v0_MV3SZ3_0 m1_499212_228525# m1_499212_228525# m1_499212_228525# m1_499212_228525#
+ VSUBS diode_nd2ps_06v0_MV3SZ3$2
Xdiode_pd2nw_06v0_5DG9HC_0 m1_499212_228525# m1_499212_228525# m1_497955_232243# m1_499212_228525#
+ m1_499212_228525# diode_pd2nw_06v0_5DG9HC$2
.ends

.subckt M a_408568_255933# a_365828_259091# a_411044_251737# a_409618_256263# a_404831_244568#
+ a_401271_243528# a_409818_256643# a_365828_265695# a_376520_259212# a_395682_259299#
+ a_411044_242557# w_364522_258756#
X0 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0.4068n ps=1.46136m w=10u l=2u
X1 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X2 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X3 a_402461_244568# a_401271_243528# a_401941_244568# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X4 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X5 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X6 a_404311_244568# a_401151_244568# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X7 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X8 a_374398_259299# a_365828_259091# a_373878_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X9 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X10 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X11 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X12 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X13 a_401151_244568# a_401151_244568# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X14 a_404041_244568# a_409618_256263# a_409618_260539# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X15 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.64p pd=17.16u as=0.1744n ps=0.65672m w=8u l=1u
X16 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X17 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X18 a_409618_256263# a_409618_260539# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X19 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X20 a_409618_256263# a_409498_256643# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X21 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X22 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X23 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X24 a_409618_256263# a_409618_260539# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X25 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X26 a_401151_244568# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X27 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X28 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X29 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X30 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X31 a_401151_244568# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X32 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X33 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X34 a_404041_244568# a_401271_243528# a_403521_244568# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X35 a_395162_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X36 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X37 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X38 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X39 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X40 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X41 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X42 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X43 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X44 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X45 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X46 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X47 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X48 a_402731_244568# a_401151_244568# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X49 a_365708_259299# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X50 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X51 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X52 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X53 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X54 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X55 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X56 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X57 a_409498_256643# a_404041_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X58 a_395682_259299# a_383940_262205# a_395162_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X59 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X60 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X61 a_409618_260539# a_404041_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X62 a_401941_244568# a_401151_244568# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X63 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X64 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X65 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X66 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X67 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X68 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X69 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X70 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X71 a_409618_260539# a_404041_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X72 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X73 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X74 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X75 a_411044_242557# a_402461_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X76 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X77 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X78 a_401151_244568# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X79 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X80 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X81 a_402461_244568# a_402461_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X82 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X83 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X84 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X85 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X86 a_404041_244568# a_409618_256263# a_409618_260539# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X87 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X88 a_404831_244568# a_401271_243528# a_404311_244568# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X89 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X90 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X91 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X92 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X93 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X94 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X95 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X96 a_401271_243528# a_401271_243528# a_401151_244568# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X97 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X98 a_403521_244568# a_401151_244568# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X99 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X100 a_365708_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X101 a_410724_251737# a_410134_251737# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X102 a_409618_256263# a_409498_256643# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X103 a_411044_251737# a_403251_244568# a_410724_251737# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X104 a_409818_256643# a_409618_256263# a_409498_256643# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X105 a_386992_259299# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X106 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X107 a_410134_251737# a_410134_251737# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X108 a_403251_244568# a_403251_244568# a_410134_251737# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X109 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X110 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X111 a_409818_256643# a_409618_256263# a_409498_256643# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X112 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X113 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X114 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X115 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X116 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X117 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X118 a_376520_259212# a_376520_259212# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.32p pd=9.16u as=0 ps=0 w=4u l=1u
X119 a_383940_262205# a_383940_262205# a_386992_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X120 a_365828_259091# a_365828_259091# a_365708_259299# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X121 a_383620_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X122 a_377450_262205# a_377450_262205# a_376520_259212# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X123 a_373878_259299# a_365708_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X124 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X125 a_409498_256643# a_404041_244568# a_376520_259212# a_376520_259212# nfet_03v3 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=1u
X126 a_401151_244568# a_365828_265695# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X127 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X128 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X129 w_364522_258756# w_364522_258756# w_364522_258756# w_364522_258756# pfet_03v3 ad=5.8p pd=21.16u as=0 ps=0 w=10u l=2u
X130 a_403251_244568# a_401271_243528# a_402731_244568# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X131 a_386992_259299# a_386992_259299# w_364522_258756# w_364522_258756# pfet_03v3 ad=6p pd=21.2u as=6p ps=21.2u w=10u l=2u
X132 a_383940_262205# a_374398_259299# a_383620_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X133 a_374398_259299# a_374398_259299# a_377450_262205# a_376520_259212# nfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
.ends

.subckt TOP CCM_OUT PU VDD VSS VIN_OUT BCM_OUT VCM_OUT VIN VBIAS EN PD
Xsc_tieh_tiel$1_0 PD PU VDD VSS sc_tieh_tiel$1
Xio_secondary_5p0$1_0 m3_419992_265695# VDD EN VSS io_secondary_5p0$1
XM_0 VSS a_499016_248165# BCM_OUT m4_400150_261569# VIN_OUT a_498947_268180# CCM_OUT
+ m3_419992_265695# VSS m4_400150_261569# VCM_OUT VDD M
D0 a_498947_268180# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D1 a_498947_268180# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D2 VSS a_499016_248165# diode_nd2ps_06v0 pj=40u area=99.99999p
X0 a_498947_268180# VIN VDD ppolyf_u r_width=40u r_length=10u
D3 a_499016_248165# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D4 a_499016_248165# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D5 VSS a_499016_248165# diode_nd2ps_06v0 pj=40u area=99.99999p
D6 a_498947_268180# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D7 VSS a_498947_268180# diode_nd2ps_06v0 pj=40u area=99.99999p
D8 a_499016_248165# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D9 a_499016_248165# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
D10 VSS a_498947_268180# diode_nd2ps_06v0 pj=40u area=99.99999p
D11 VSS a_499016_248165# diode_nd2ps_06v0 pj=40u area=99.99999p
D12 VSS a_498947_268180# diode_nd2ps_06v0 pj=40u area=99.99999p
D13 a_498947_268180# VDD diode_pd2nw_06v0 pj=40u area=99.99999p
X1 a_499016_248165# VBIAS VDD ppolyf_u r_width=40u r_length=10u
D14 VSS a_499016_248165# diode_nd2ps_06v0 pj=40u area=99.99999p
D15 VSS a_498947_268180# diode_nd2ps_06v0 pj=40u area=99.99999p
.ends

