| units: 0.5 tech: gf180mcuD format: MIT
x a_n2573_n881# VDD a_n2573_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=1677 y=1625 pfet_03v3
x VIN a_n2573_n881# VIN VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=1677 y=-880 pfet_03v3
x VIN a_n2573_n881# VIN VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=2857 y=-880 pfet_03v3
x a_n2573_n881# VDD a_n2573_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=2857 y=1625 pfet_03v3
x VIN a_n2573_n881# VIN VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=-1862 y=-880 pfet_03v3
x a_n2573_n881# VDD a_n2573_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=-1862 y=1625 pfet_03v3
x a_n2573_n881# VDD a_n2573_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=1087 y=1625 pfet_03v3
x VIN a_n2573_n881# VIN VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=1087 y=-880 pfet_03v3
x VIN a_n2573_n881# VIN VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=2267 y=-880 pfet_03v3
x a_n2573_n881# VDD a_n2573_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=2267 y=1625 pfet_03v3
x VIN a_n2573_n881# VIN VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=-1272 y=-880 pfet_03v3
x a_n2573_n881# VDD a_n2573_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=-2452 y=1625 pfet_03v3
x a_n2573_n881# VDD a_n2573_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=-1272 y=1625 pfet_03v3
x VIN a_n2573_n881# VIN VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=-2452 y=-880 pfet_03v3
x a_n2573_n881# VDD a_n2573_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=-92 y=1625 pfet_03v3
x VIN a_n2573_n881# VIN VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=-92 y=-880 pfet_03v3
x VDD VDD VDD VDD d=185600,3432 l=200 w=1600 x=-3060 y=1625 pfet_03v3
x a_n2573_n881# VDD a_n2573_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=-682 y=1625 pfet_03v3
x a_n2573_n881# VDD a_n2573_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=497 y=1625 pfet_03v3
x VDD VDD VDD VDD d=185600,3432 l=200 w=1600 x=-3060 y=-880 pfet_03v3
x VIN a_n2573_n881# VIN VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=-682 y=-880 pfet_03v3
x VIN a_n2573_n881# VIN VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=497 y=-880 pfet_03v3
x VIN a_3597_n881# VOUT VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=3717 y=-880 pfet_03v3
x a_n2573_n881# VDD a_3597_n881# VDD s=192000,3440 d=192000,3440 l=200 w=1600 x=3717 y=1625 pfet_03v3
x VDD VDD VDD VDD d=185600,3432 l=200 w=1600 x=4325 y=-880 pfet_03v3
x VDD VDD VDD VDD d=185600,3432 l=200 w=1600 x=4325 y=1625 pfet_03v3
C a_3597_n881# VIN 0.7
C VDD a_n2573_n881# 38.2
C VDD VOUT 1.2
C VDD VIN 10.8
C a_n2573_n881# VOUT 0.0
C a_n2573_n881# VIN 26.2
C VIN VOUT 0.3
C VDD a_3597_n881# 2.9
C a_n2573_n881# a_3597_n881# 0.7
C a_3597_n881# VOUT 1.0
C VOUT0 0.3
R VOUT 99
C VIN0 1.5
R VIN 2035
C VDD0 142.3
R VDD 6445
C a_3597_n881#0 0.3
R a_3597_n881# 212
C a_n2573_n881#0 1.5
R a_n2573_n881# 3161
