** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/dc_lv_nmos.sch
**.subckt dc_lv_nmos
Vgs G GND 1.2
Vds D GND 1.5
Vd D net1 0
.save i(vd)
XM1 net1 G GND GND sg13_lv_nmos w=1.0u l=2.0u ng=1 m=1
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.include dc_lv_nmos.save
.param temp=27
.control
save all
op
write dc_lv_nmos.raw
set appendwrite
*dc Vds 0 1.2 0.01 Vgs 0.3 1.0 0.1
dc Vgs 0 0.5 0.05
write dc_lv_nmos.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
