** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/neuron_buff_test.sch
**.subckt neuron_buff_test
XM3 vmem VLK GND GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=1
XM1 GND VTHR vn1 VDD sg13_lv_pmos w=1.2u l=0.75u ng=1 m=1
XM4 vmem vmem vn1 VDD sg13_lv_pmos w=1.2u l=0.75u ng=1 m=1
Vdd1 VDD GND 1.8
XM24 VREF VREF GND GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=1
IVREF VDD VREF 700nA
XM5 vmem RST GND GND sg13_lv_nmos w=1.2u l=0.28u ng=1 m=1
XM6 net2 net1 VDD VDD sg13_lv_pmos w=2.4u l=3.0u ng=1 m=1
XM8 vmem REQ net2 VDD sg13_lv_pmos w=2.4u l=0.28u ng=1 m=1
XM9 net1 net1 VDD VDD sg13_lv_pmos w=2.4u l=3.0u ng=1 m=1
XM10 REQ vmem net1 VDD sg13_lv_pmos w=2.4u l=0.28u ng=1 m=1
XM11 REQ vmem net3 GND sg13_lv_nmos w=1.2u l=0.28u ng=1 m=1
XM25 net3 net3 GND GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=1
XM26 net4 REQ net6 VDD sg13_lv_pmos w=2.4u l=0.28u ng=1 m=1
XM27 net4 REQ net5 GND sg13_lv_nmos w=1.2u l=0.28u ng=1 m=1
XM28 net5 VREF GND GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=1
XM29 net6 net6 net7 VDD sg13_lv_pmos w=2.4u l=3.0u ng=1 m=1
XM30 net7 REQ VDD VDD sg13_lv_pmos w=2.4u l=0.28u ng=1 m=1
xinv2 VDD net11 net12 GND inv
* noconn OUT
XM2 VTHR VTHR GND GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=1
ITHR VDD VTHR 300n
XM7 net8 net4 net9 VDD sg13_lv_pmos w=2.4u l=0.28u ng=1 m=1
XM12 net8 net4 GND GND sg13_lv_nmos w=1.2u l=0.28u ng=1 m=1
XM14 net9 net9 VDD VDD sg13_lv_pmos w=2.4u l=3.0u ng=1 m=1
XM13 RST net8 net10 VDD sg13_lv_pmos w=2.4u l=0.28u ng=1 m=1
XM15 RST net8 GND GND sg13_lv_nmos w=1.2u l=0.28u ng=1 m=1
XM16 net10 net10 VDD VDD sg13_lv_pmos w=2.4u l=3.0u ng=1 m=1
XM17 GND vmem GND GND sg13_lv_pmos w=5.0u l=10.0u ng=6 m=10
XM18 GND RST GND GND sg13_lv_pmos w=5.0u l=10.0u ng=6 m=10
xinv1 VDD REQ net11 GND inv
xinv3 net21 net12 OUT GND inv
xinv4 VDD net11 net12 GND inv
xinv5 VDD net12 OUT GND inv
Ven6 DB0 GND 1.8
Ven7 DB1 GND 0
Ven8 DB2 GND 0
Ven9 DB3 GND 0
x2 DB0 DB1 DB2 DB3 VDD GND CSen2 net19 trimmer
Ven5 CSen2 GND 1.8
XM35 net13 net13 net14 GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=10
XM36 net16 net13 net15 GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=1
XM37 net14 net14 GND GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=10
XM38 net15 net14 GND GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=1
XM39 net16 net16 net17 VDD sg13_lv_pmos w=2.4u l=3.0u ng=1 m=10
XM40 net20 net16 net18 VDD sg13_lv_pmos w=2.4u l=3.0u ng=1 m=1
XM41 net17 net17 VDD VDD sg13_lv_pmos w=2.4u l=3.0u ng=1 m=10
XM42 net18 net17 VDD VDD sg13_lv_pmos w=2.4u l=3.0u ng=1 m=1
XM23 VLK VLK GND GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=1
IVREF1 VDD vn1 30nA
Vmeas net19 net13 0
.save i(vmeas)
Vmeas1 net20 VLK 0
.save i(vmeas1)
XM33 ob1 ob1 GND GND sg13_lv_nmos w=1.2u l=3.0u ng=1 m=1
ILK VDD ob1 3nA
* noconn ob1
**** begin user architecture code

.include diodes.lib
.include sg13g2_bondpad.lib



.options savecurrents
.include neuron_buff_test.save
.param temp=27
.control
set wr_singlescale
set noaskquit
*set appendwrite
set hcopypscolor=1

*Save node voltages and device currents if desired
save all

*Baseline operating point at current deck values
op
write tran_neuron.raw

alter Ven dc 1.8
alter ven6 dc 1.8
alter ven7 dc 0.0
alter ven8 dc 0.0
alter ven9 dc 0.0

tran 1u 100u
write tran_neuron.raw
*Example plots (uncomment inside ngspice if you want autoplots)
plot vmem vn1 Vthr Vlk
plot vmem out
plot vmeas1#branch vmeas2#branch vmeas3#branch vmeas4#branch
*quit
.endc





.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ


**** end user architecture code
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/inv.sym
** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/inv.sch
.subckt inv VDD in out VSS
*.iopin VDD
*.ipin in
*.iopin VSS
*.opin out
XM1 out in VSS VSS sg13_lv_nmos w=1.2u l=0.28u ng=1 m=1
XM2 out in VDD VDD sg13_lv_pmos w=2.4u l=0.28u ng=1 m=1
.ends


* expanding   symbol:  trimmer.sym # of pins=8
** sym_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/trimmer.sym
** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/trimmer.sch
.subckt trimmer D0 D1 D2 D3 VDD VSS en out
*.ipin en
*.ipin D0
*.ipin D1
*.ipin D2
*.ipin D3
*.opin out
*.iopin VDD
*.iopin VSS
XMP1 net1 net1 net12 VDD sg13_lv_pmos w=0.28u l=8.0u ng=1 m=1
XMP2 vstart vstart net1 VDD sg13_lv_pmos w=0.28u l=8.0u ng=1 m=1
XMN2 net3 vstart GND GND sg13_lv_nmos w=0.28u l=8.0u ng=1 m=1
XMN1 vstart vstart GND GND sg13_lv_nmos w=0.28u l=8.0u ng=1 m=1
XMP3 net2 vbp net11 VDD sg13_lv_pmos w=2.0u l=2.0u ng=2 m=1
XMP4 net3 vbp_casc net2 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP5 net4 vbp net10 VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=2
XMP6 net6 vbp_casc net4 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP7 net5 vbp net9 VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=2
XMP8 vbp vbp_casc net5 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP9 net6 net3 VDD VDD sg13_lv_pmos w=0.28u l=8.0u ng=1 m=1
XMN3 net6 net6 GND GND sg13_lv_nmos w=2.0u l=2.0u ng=1 m=1
XMN4 vbp_casc net6 net7 GND sg13_lv_nmos w=2.0u l=2.0u ng=1 m=4
XR1 vbp_casc vbp sub! rppd w=0.5e-6 l=389e-6 m=1 b=0
XR2 GND net7 sub! rhigh w=0.5e-6 l=152.5e-6 m=1 b=0
XMP10 net13 vbp net14 VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=2
XMP11 out vbp_casc net13 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP16 vbp_casc enMon VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=1
XMP17 net9 net8 VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP18 net10 net8 VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP19 net12 net8 VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=1
XMP20 net11 net8 VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=1
XMN5 vstart net8 GND GND sg13_lv_nmos w=2u l=0.28u ng=1 m=1
XMN6 net6 net8 GND GND sg13_lv_nmos w=2u l=0.28u ng=1 m=1
xinv2 VDD net8 enMon GND inv
XMP12 net14 net15 VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP13 net16 vbp net17 VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=4
XMP14 out vbp_casc net16 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=4
XMP15 net17 net18 VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP21 net19 vbp net20 VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=8
XMP22 out vbp_casc net19 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=8
XMP23 net20 net21 VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
XMP24 net22 vbp net23 VDD sg13_lv_pmos w=2.0u l=2.0u ng=1 m=16
XMP25 out vbp_casc net22 VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=16
XMP26 net23 net24 VDD VDD sg13_lv_pmos w=2.0u l=0.28u ng=1 m=2
xinv6 VDD en net8 GND inv
xinv3 VDD D0 net15 GND inv
xinv7 VDD D1 net18 GND inv
xinv8 VDD D2 net21 GND inv
xinv9 VDD D3 net24 GND inv
.ends

.GLOBAL GND
.GLOBAL VDD
.end
