| units: 0.5 tech: gf180mcuD format: MIT
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=-1002 y=-584 nfet_03v3
x VIN a_75_1553# VOUT VSS s=96000,1840 d=96000,1840 l=200 w=800 x=195 y=1553 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=803 y=-584 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=-1002 y=1553 nfet_03v3
x a_n515_1553# VSS a_n515_1553# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=-394 y=-584 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=803 y=1553 nfet_03v3
x a_n515_1553# VSS a_75_1553# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=195 y=-584 nfet_03v3
x VIN a_n515_1553# VIN VSS s=96000,1840 d=96000,1840 l=200 w=800 x=-394 y=1553 nfet_03v3
C VIN a_n515_1553# 1.8
C a_75_1553# a_n515_1553# 0.4
C VIN VOUT 0.2
C a_75_1553# VOUT 1.2
C a_75_1553# VIN 1.5
C VOUT a_n515_1553# 0.1
C VOUT0 1.7
R VOUT 47
C VIN0 2.7
R VIN 159
R VSS 2236
C a_75_1553#0 2.9
R a_75_1553# 107
C a_n515_1553#0 6.5
R a_n515_1553# 219
