| units: 0.5 tech: gf180mcuD format: MIT
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2587 y=-1499 pfet_03v3
x VIN a_n1110_n1500# VOUT_VCM VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-989 y=-1499 pfet_03v3
x EN VDD a_n1900_n1500# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=195 y=9300 pfet_03v3
x VIN a_1260_n1500# VOUT_VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=1380 y=-1499 pfet_03v3
x a_n1900_n1500# VDD a_n320_n1500# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-199 y=3848 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=2188 y=3848 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2192 y=9300 pfet_03v3
x EN VDD a_n1900_n1500# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-594 y=9300 pfet_03v3
x VIN a_n320_n1500# VOUT_BCM VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-199 y=-1499 pfet_03v3
x EN VDD a_n1900_n1500# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=985 y=9300 pfet_03v3
x VIN a_n1900_n1500# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1779 y=-1499 pfet_03v3
x a_n1900_n1500# VDD a_n1110_n1500# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-989 y=3848 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2587 y=3848 pfet_03v3
x a_n1900_n1500# VDD a_470_n1500# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=590 y=3848 pfet_03v3
x EN VDD a_n1900_n1500# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1384 y=9300 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1793 y=9300 pfet_03v3
x VIN a_470_n1500# VOUT_CCM VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=590 y=-1499 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=2188 y=-1499 pfet_03v3
x a_n1900_n1500# VDD a_n1900_n1500# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1779 y=3848 pfet_03v3
x a_n1900_n1500# VDD a_1260_n1500# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=1380 y=3848 pfet_03v3
C a_n320_n1500# a_1260_n1500# 0.3
C VOUT_VIN a_n1900_n1500# 1.0
C VOUT_VIN VIN 0.5
C VDD a_470_n1500# 7.5
C VOUT_CCM a_1260_n1500# 2.3
C a_n1900_n1500# VOUT_VCM 0.1
C VOUT_BCM a_n1900_n1500# 0.1
C VIN VOUT_VCM 0.6
C VOUT_BCM VIN 0.6
C a_n320_n1500# VOUT_VIN 0.1
C EN a_n1110_n1500# 0.0
C VDD a_n1900_n1500# 44.9
C a_n320_n1500# VOUT_VCM 2.3
C VOUT_CCM VOUT_VIN 0.3
C VDD VIN 14.5
C VOUT_BCM a_n320_n1500# 2.4
C VOUT_CCM VOUT_VCM 0.1
C VOUT_BCM VOUT_CCM 0.3
C a_1260_n1500# a_n1110_n1500# 0.3
C VDD a_n320_n1500# 7.4
C a_470_n1500# a_n1900_n1500# 1.5
C a_470_n1500# VIN 0.6
C VDD VOUT_CCM 1.1
C VOUT_VIN a_n1110_n1500# 0.1
C a_n320_n1500# a_470_n1500# 0.8
C VOUT_VCM a_n1110_n1500# 2.4
C VOUT_BCM a_n1110_n1500# 0.2
C a_1260_n1500# EN 0.3
C a_n1900_n1500# VIN 3.4
C VOUT_CCM a_470_n1500# 2.4
C VDD a_n1110_n1500# 7.4
C a_n320_n1500# a_n1900_n1500# 1.5
C a_n320_n1500# VIN 0.6
C VOUT_CCM a_n1900_n1500# 0.1
C VOUT_CCM VIN 0.6
C a_470_n1500# a_n1110_n1500# 0.3
C VOUT_VIN a_1260_n1500# 2.4
C a_n320_n1500# VOUT_CCM 0.2
C VDD EN 11.1
C a_1260_n1500# VOUT_VCM 0.1
C VOUT_BCM a_1260_n1500# 0.1
C a_n1900_n1500# a_n1110_n1500# 1.8
C VIN a_n1110_n1500# 2.9
C VDD a_1260_n1500# 6.4
C a_470_n1500# EN 0.0
C VOUT_VIN VOUT_VCM 0.1
C VOUT_BCM VOUT_VIN 0.1
C a_n320_n1500# a_n1110_n1500# 0.8
C VOUT_BCM VOUT_VCM 0.3
C VOUT_CCM a_n1110_n1500# 0.2
C VDD VOUT_VIN 2.2
C a_470_n1500# a_1260_n1500# 0.8
C EN a_n1900_n1500# 2.2
C VDD VOUT_VCM 1.2
C VDD VOUT_BCM 1.1
C a_n320_n1500# EN 0.0
C a_470_n1500# VOUT_VIN 0.1
C a_1260_n1500# a_n1900_n1500# 2.4
C a_1260_n1500# VIN 0.6
C a_470_n1500# VOUT_VCM 0.1
C VOUT_BCM a_470_n1500# 2.3
C VOUT_VIN0 0.4
R VOUT_VIN 128
C VOUT_CCM0 0.2
R VOUT_CCM 128
C VOUT_BCM0 0.2
R VOUT_BCM 128
C VOUT_VCM0 0.3
R VOUT_VCM 128
C VIN0 2.5
R VIN 515
C EN0 1.8
R EN 289
C VDD0 304.6
R VDD 9768
C a_1260_n1500#0 0.2
R a_1260_n1500# 272
C a_470_n1500#0 0.0
R a_470_n1500# 272
C a_n320_n1500#0 0.0
R a_n320_n1500# 272
C a_n1110_n1500#0 0.0
R a_n1110_n1500# 272
C a_n1900_n1500#0 3.2
R a_n1900_n1500# 1220
