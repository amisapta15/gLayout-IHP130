** sch_path: /foss/designs/gLayout-IHP130/blocks/composite/dpi_adexp_neuron/design_data/xschem/sbcmN.sch
**.subckt sbcmN VDD GND IREF ICOPY
*.iopin VDD
*.iopin GND
*.iopin IREF
*.iopin ICOPY
XM6 net2 net1 VDD VDD sg13_lv_pmos w=15.0u l=0.5u ng=5 m=1
XM9 net3 net1 VDD VDD sg13_lv_pmos w=15.0u l=0.5u ng=5 m=10
XM1 ICOPY IREF net2 VDD sg13_lv_pmos w=15.0u l=0.5u ng=5 m=1
XM2 net1 IREF net3 VDD sg13_lv_pmos w=15.0u l=0.5u ng=5 m=10
XM23 net1 VDD IREF GND sg13_lv_nmos w=21.0u l=0.5u ng=7 m=10
XM3 net4 net4 net5 GND sg13_lv_nmos w=8.0u l=0.5u ng=1 m=10
XM4 net7 net4 net6 GND sg13_lv_nmos w=8.0u l=0.5u ng=1 m=1
XM5 net5 net5 GND GND sg13_lv_nmos w=8.0u l=0.5u ng=1 m=10
XM7 net6 net5 GND GND sg13_lv_nmos w=8.0u l=0.5u ng=1 m=1
I0 VDD net4 300n
V1 net7 GND 0
**** begin user architecture code


.include sbcmN.save
.option savecurrent
.param temp=127
.control
save all
op
write sbcmN.raw
*tran 1n 5u
dc V1 0 1.8 0.1
write sbcmN.raw
plot -i(V1)
.endc





.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ


**** end user architecture code
**.ends
.end
