magic
tech gf180mcuD
magscale 1 10
timestamp 1757928106
<< nwell >>
rect -4460 -1160 4460 1160
<< pwell >>
rect -4622 1160 4622 1322
rect -4622 -1160 -4460 1160
rect 4460 -1160 4622 1160
rect -4622 -1322 4622 -1160
<< psubdiff >>
rect -4598 1285 4598 1298
rect -4598 1239 -4482 1285
rect 4482 1239 4598 1285
rect -4598 1226 4598 1239
rect -4598 1182 -4526 1226
rect -4598 -1182 -4585 1182
rect -4539 -1182 -4526 1182
rect 4526 1182 4598 1226
rect -4598 -1226 -4526 -1182
rect 4526 -1182 4539 1182
rect 4585 -1182 4598 1182
rect 4526 -1226 4598 -1182
rect -4598 -1239 4598 -1226
rect -4598 -1285 -4482 -1239
rect 4482 -1285 4598 -1239
rect -4598 -1298 4598 -1285
<< nsubdiff >>
rect -4436 1123 4436 1136
rect -4436 1073 -4316 1123
rect -2284 1073 -2116 1123
rect -84 1073 84 1123
rect 2116 1073 2284 1123
rect 4316 1073 4436 1123
rect -4436 1060 4436 1073
rect -4436 1016 -4360 1060
rect -4436 -1016 -4423 1016
rect -4373 -1016 -4360 1016
rect -2240 1016 -2160 1060
rect -4436 -1060 -4360 -1016
rect -2240 -1016 -2227 1016
rect -2173 -1016 -2160 1016
rect -40 1016 40 1060
rect -2240 -1060 -2160 -1016
rect -40 -1016 -27 1016
rect 27 -1016 40 1016
rect 2160 1016 2240 1060
rect -40 -1060 40 -1016
rect 2160 -1016 2173 1016
rect 2227 -1016 2240 1016
rect 4360 1016 4436 1060
rect 2160 -1060 2240 -1016
rect 4360 -1016 4373 1016
rect 4423 -1016 4436 1016
rect 4360 -1060 4436 -1016
rect -4436 -1073 4436 -1060
rect -4436 -1123 -4316 -1073
rect -2284 -1123 -2116 -1073
rect -84 -1123 84 -1073
rect 2116 -1123 2284 -1073
rect 4316 -1123 4436 -1073
rect -4436 -1136 4436 -1123
<< psubdiffcont >>
rect -4482 1239 4482 1285
rect -4585 -1182 -4539 1182
rect 4539 -1182 4585 1182
rect -4482 -1285 4482 -1239
<< nsubdiffcont >>
rect -4316 1073 -2284 1123
rect -2116 1073 -84 1123
rect 84 1073 2116 1123
rect 2284 1073 4316 1123
rect -4423 -1016 -4373 1016
rect -2227 -1016 -2173 1016
rect -27 -1016 27 1016
rect 2173 -1016 2227 1016
rect 4373 -1016 4423 1016
rect -4316 -1123 -2284 -1073
rect -2116 -1123 -84 -1073
rect 84 -1123 2116 -1073
rect 2284 -1123 4316 -1073
<< pdiode >>
rect -4300 987 -2300 1000
rect -4300 -987 -4287 987
rect -2313 -987 -2300 987
rect -4300 -1000 -2300 -987
rect -2100 987 -100 1000
rect -2100 -987 -2087 987
rect -113 -987 -100 987
rect -2100 -1000 -100 -987
rect 100 987 2100 1000
rect 100 -987 113 987
rect 2087 -987 2100 987
rect 100 -1000 2100 -987
rect 2300 987 4300 1000
rect 2300 -987 2313 987
rect 4287 -987 4300 987
rect 2300 -1000 4300 -987
<< pdiodec >>
rect -4287 -987 -2313 987
rect -2087 -987 -113 987
rect 113 -987 2087 987
rect 2313 -987 4287 987
<< metal1 >>
rect -4585 1239 -4482 1285
rect 4482 1239 4585 1285
rect -4585 1182 -4539 1239
rect 4539 1182 4585 1239
rect -4423 1073 -4316 1123
rect -2284 1073 -2116 1123
rect -84 1073 84 1123
rect 2116 1073 2284 1123
rect 4316 1073 4423 1123
rect -4423 1016 -4373 1073
rect -2227 1016 -2173 1073
rect -4298 -987 -4287 987
rect -2313 -987 -2302 987
rect -4423 -1073 -4373 -1016
rect -27 1016 27 1073
rect -2098 -987 -2087 987
rect -113 -987 -102 987
rect -2227 -1073 -2173 -1016
rect 2173 1016 2227 1073
rect 102 -987 113 987
rect 2087 -987 2098 987
rect -27 -1073 27 -1016
rect 4373 1016 4423 1073
rect 2302 -987 2313 987
rect 4287 -987 4298 987
rect 2173 -1073 2227 -1016
rect 4373 -1073 4423 -1016
rect -4423 -1123 -4316 -1073
rect -2284 -1123 -2116 -1073
rect -84 -1123 84 -1073
rect 2116 -1123 2284 -1073
rect 4316 -1123 4423 -1073
rect -4585 -1239 -4539 -1182
rect 4539 -1239 4585 -1182
rect -4585 -1285 -4482 -1239
rect 4482 -1285 4585 -1239
<< properties >>
string diode_pd2nw_03v3_5DG9GA parameters
string FIXED_BBOX 2202 -1098 4398 1098
string gencell diode_pd2nw_03v3
string library gf180mcu
string parameters w 10 l 10 area 100.0 peri 40.0 nx 4 ny 1 dummy 0 lmin 0.45 wmin 0.45 class diode elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 1 full_metal 1 compatible {diode_pd2nw_03v3 diode_pd2nw_06v0}
<< end >>
