* NGSPICE file created from M.ext - technology: sky130A

.subckt M VIN VSS VDD VOUT_VIN VOUT_RCCM VOUT_SBCM VOUT_VCM VAUX EN
X0 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X1 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=115.44 ps=634.90002 w=4 l=1
X2 a_n17107_9910# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X3 a_200_n5640# a_200_n5640# a_6260_503# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X4 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X5 VOUT_RCCM a_5835_4440# a_5757_4829# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X6 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=81.9078 ps=436.42001 w=10 l=2
X7 a_n32245_7124# EN w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X8 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X9 a_6722_503# a_6260_503# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X10 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X11 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X12 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X13 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X14 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X15 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X16 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X17 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X18 a_5835_4440# a_5757_4829# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X19 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X20 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X21 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=0 ps=0 w=10.005 l=2
X22 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=187.2 ps=997.44 w=10 l=2
X23 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=0 ps=0 w=10.005 l=2
X24 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X25 a_n1602_n5640# EN w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X26 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X27 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X28 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X29 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X30 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X31 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X32 a_5835_8163# a_862_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X33 a_n1602_n5640# EN w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X34 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X35 VOUT_VCM a_n462_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X36 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X37 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X38 a_5757_4829# a_862_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X39 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X40 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X41 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X42 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X43 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X44 a_5835_4440# a_5835_8163# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X45 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X46 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X47 a_n278_n5640# a_n1602_n5640# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X48 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X49 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X50 a_1046_n5640# a_n1602_n5640# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X51 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X52 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X53 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X54 a_200_n5640# a_n1524_n6691# a_n278_n5640# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=3.90195 ps=20.79 w=10.005 l=2
X55 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X56 a_384_n5640# a_n1602_n5640# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X57 a_862_n5640# a_5835_4440# a_5835_8163# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X58 a_6260_503# a_6260_503# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X59 a_n6641_7124# a_n16829_9910# a_n7119_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X60 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X61 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X62 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X63 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X64 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X65 a_n1602_n5640# EN w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X66 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X67 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X68 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X69 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X70 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X71 VOUT_VIN a_n1524_n6691# a_1046_n5640# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=3.90195 ps=20.79 w=10.005 l=2
X72 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X73 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X74 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X75 a_n24817_7124# VAUX a_n25295_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X76 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X77 VOUT_RCCM a_5835_4440# a_5757_4829# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X78 a_n462_n5640# a_n462_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X79 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X80 a_5835_4440# a_5757_4829# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X81 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X82 a_n1524_n6691# a_n1524_n6691# a_n1602_n5640# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=3.90195 ps=20.79 w=10.005 l=2
X83 a_n940_n5640# a_n1602_n5640# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X84 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X85 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X86 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X87 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X88 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X89 a_n1602_n5640# a_n1602_n5640# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X90 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X91 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X92 a_n16829_9910# a_n24817_7124# a_n17107_9910# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X93 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X94 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X95 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X96 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X97 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X98 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X99 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X100 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X101 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X102 a_5835_8163# a_862_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X103 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X104 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X105 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X106 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X107 a_5757_4829# a_862_n5640# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X108 a_n32245_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X109 a_n7119_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X110 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X111 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X112 a_n22057_9909# a_n22057_9909# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X113 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X114 a_n24817_7124# a_n24817_7124# a_n22057_9909# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=3.12 ps=16.78 w=8 l=1
X115 VOUT_SBCM a_200_n5640# a_6722_503# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X116 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=1
X117 w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X118 a_5835_4440# a_5835_8163# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X119 a_n462_n5640# a_n1524_n6691# a_n940_n5640# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=3.90195 ps=20.79 w=10.005 l=2
X120 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X121 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X122 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X123 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X124 a_n25295_7124# a_n32245_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X125 a_n14069_7124# a_n14069_7124# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X126 a_n22897_6995# a_n22897_6995# a_n22897_6995# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X127 VAUX VAUX a_n32245_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X128 a_862_n5640# a_5835_4440# a_5835_8163# a_n22897_6995# sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=1
X129 w_n33347_6533# w_n33347_6533# w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=2
X130 a_862_n5640# a_n1524_n6691# a_384_n5640# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.90195 pd=20.79 as=3.90195 ps=20.79 w=10.005 l=2
X131 a_n14069_7124# EN w_n33347_6533# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X132 a_n1602_n5640# EN w_n2704_n7119# w_n2704_n7119# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
X133 a_n16829_9910# a_n16829_9910# a_n14069_7124# w_n33347_6533# sky130_fd_pr__pfet_01v8 ad=3.9 pd=20.78 as=3.9 ps=20.78 w=10 l=2
.ends

