* NGSPICE file created from BB.ext - technology: gf180mcuD

.subckt BB VIN VDD VOUT
X0 a_n2573_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X1 VIN VIN a_n2573_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X2 VIN VIN a_n2573_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X3 a_n2573_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X4 VIN VIN a_n2573_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X5 a_n2573_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X6 a_n2573_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X7 VIN VIN a_n2573_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X8 VIN VIN a_n2573_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X9 a_n2573_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X10 VIN VIN a_n2573_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X11 a_n2573_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X12 a_n2573_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X13 VIN VIN a_n2573_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X14 a_n2573_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X15 VIN VIN a_n2573_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X16 VDD VDD VDD VDD pfet_03v3 ad=4.64p pd=17.16u as=89.92p ps=0.32648m w=8u l=1u
X17 a_n2573_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X18 a_n2573_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X19 VDD VDD VDD VDD pfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X20 VIN VIN a_n2573_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X21 VIN VIN a_n2573_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X22 VOUT VIN a_3597_n881# VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X23 a_3597_n881# a_n2573_n881# VDD VDD pfet_03v3 ad=4.8p pd=17.2u as=4.8p ps=17.2u w=8u l=1u
X24 VDD VDD VDD VDD pfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
X25 VDD VDD VDD VDD pfet_03v3 ad=4.64p pd=17.16u as=0 ps=0 w=8u l=1u
.ends

