| units: 0.5 tech: gf180mcuD format: MIT
x a_5777_8307# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=5777 y=8687 nfet_03v3
x a_5777_8307# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6957 y=8687 nfet_03v3
x a_5657_4411# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6367 y=4411 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5805 y=-7718 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2192 y=-1233 pfet_03v3
x a_n1505_n5930# VDD a_n715_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-594 y=-1233 pfet_03v3
x a_5657_4411# VSS VAUX VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7547 y=4411 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=7611 y=-1654 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1793 y=-1233 pfet_03v3
x VIN a_n715_n5930# a_n195_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-594 y=-5929 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5169 y=4411 nfet_03v3
x a_n1505_n5930# VDD a_75_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=195 y=-1233 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-2192 y=-5929 pfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1793 y=-5929 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=7611 y=-7718 nfet_03v3
x VAUX a_5777_8307# a_1385_n5930# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6367 y=8687 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8155 y=4411 nfet_03v3
x a_595_n5930# a_6293_483# a_595_n5930# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6413 y=483 nfet_03v3
x EN VDD a_n1505_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-199 y=3567 pfet_03v3
x VIN a_75_n5930# a_595_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=195 y=-5929 pfet_03v3
x VAUX a_5777_8307# a_1385_n5930# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7547 y=8687 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5169 y=8687 nfet_03v3
x a_6293_483# VSS a_6883_483# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7003 y=-1654 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8155 y=8687 nfet_03v3
x a_1385_n5930# VSS a_5777_8307# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=5777 y=6549 nfet_03v3
x a_1385_n5930# VSS a_5777_8307# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6957 y=6549 nfet_03v3
x a_n195_n5930# VSS VOUT_VCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7003 y=-7718 nfet_03v3
x a_595_n5930# a_6883_483# VOUT_SBCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7003 y=483 nfet_03v3
x a_1385_n5930# VSS a_5657_4411# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6367 y=6549 nfet_03v3
x a_1385_n5930# VSS a_5657_4411# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=7547 y=6549 nfet_03v3
x EN VDD a_n1505_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-989 y=3567 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5169 y=6549 nfet_03v3
x a_n1505_n5930# VDD a_n1505_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1384 y=-1233 pfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=8155 y=6549 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=1398 y=3567 pfet_03v3
x VIN a_n1505_n5930# VIN VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=-1384 y=-5929 pfet_03v3
x EN VDD a_n1505_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=590 y=3567 pfet_03v3
x a_n1505_n5930# VDD a_865_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=985 y=-1233 pfet_03v3
x a_6293_483# VSS a_6293_483# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6413 y=-1654 nfet_03v3
x VIN a_865_n5930# a_1385_n5930# VDD s=240000,4240 d=240000,4240 l=400 w=2000 x=985 y=-5929 pfet_03v3
x a_n195_n5930# VSS a_n195_n5930# VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6413 y=-7718 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5805 y=483 nfet_03v3
x VAUX a_5657_4411# VOUT_RCCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=5777 y=4411 nfet_03v3
x VDD VDD VDD VDD d=232000,4232 l=400 w=2000 x=-1797 y=3567 pfet_03v3
x VAUX a_5657_4411# VOUT_RCCM VSS s=96000,1840 d=96000,1840 l=200 w=800 x=6957 y=4411 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=7611 y=483 nfet_03v3
x VSS VSS VSS VSS d=92800,1832 l=200 w=800 x=5805 y=-1654 nfet_03v3
C a_n195_n5930# a_595_n5930# 0.5
C VOUT_RCCM a_5777_8307# 0.0
C VIN VDD 10.3
C a_n1505_n5930# VDD 31.5
C a_75_n5930# a_1385_n5930# 0.1
C a_n715_n5930# VDD 6.3
C a_5657_4411# a_1385_n5930# 0.9
C a_865_n5930# a_595_n5930# 2.0
C a_n195_n5930# VIN 0.6
C a_n1505_n5930# a_n195_n5930# 0.1
C a_n715_n5930# a_n195_n5930# 2.0
C a_n1505_n5930# EN 1.6
C VDD a_1385_n5930# 2.6
C a_6293_483# a_595_n5930# 1.9
C a_5777_8307# VAUX 3.6
C a_n715_n5930# EN 0.0
C a_75_n5930# VDD 6.4
C a_865_n5930# VIN 0.6
C a_865_n5930# a_n1505_n5930# 2.2
C a_865_n5930# a_n715_n5930# 0.3
C a_n195_n5930# a_1385_n5930# 0.1
C VOUT_RCCM VAUX 0.6
C a_75_n5930# a_n195_n5930# 2.0
C a_5777_8307# a_1385_n5930# 3.0
C a_6883_483# VOUT_SBCM 1.2
C VOUT_VCM a_n195_n5930# 0.2
C VIN a_595_n5930# 0.6
C a_n1505_n5930# a_595_n5930# 0.1
C a_75_n5930# EN 0.0
C a_n715_n5930# a_595_n5930# 0.2
C a_865_n5930# a_1385_n5930# 2.0
C a_5777_8307# a_5657_4411# 0.4
C a_865_n5930# a_75_n5930# 0.7
C VOUT_RCCM a_1385_n5930# 0.0
C a_n195_n5930# VDD 1.1
C a_n1505_n5930# VIN 3.0
C VDD EN 7.3
C a_595_n5930# a_1385_n5930# 0.4
C a_n715_n5930# VIN 2.6
C a_n1505_n5930# a_n715_n5930# 1.7
C VOUT_RCCM a_5657_4411# 2.2
C a_75_n5930# a_595_n5930# 2.0
C a_6883_483# a_6293_483# 0.4
C a_865_n5930# VDD 5.4
C a_6883_483# a_595_n5930# 1.5
C VIN a_1385_n5930# 0.6
C a_n1505_n5930# a_1385_n5930# 0.8
C VAUX a_1385_n5930# 1.7
C a_n715_n5930# a_1385_n5930# 0.1
C a_75_n5930# VIN 0.6
C a_865_n5930# a_n195_n5930# 0.1
C a_n1505_n5930# a_75_n5930# 1.4
C VDD a_595_n5930# 1.0
C a_5657_4411# VAUX 3.3
C VOUT_SBCM a_6293_483# 0.1
C a_n715_n5930# a_75_n5930# 0.8
C a_865_n5930# EN 0.2
C VOUT_SBCM a_595_n5930# 0.2
C VOUT_VCM0 3.0
R VOUT_VCM 47
C VOUT_SBCM0 1.7
R VOUT_SBCM 47
C VOUT_RCCM0 3.1
R VOUT_RCCM 107
C VAUX0 16.1
R VAUX 476
C VIN0 2.1
R VIN 414
C EN0 1.4
R EN 198
C VDD0 234.0
R VDD 9009
R VSS 7334
C a_6883_483#0 2.9
R a_6883_483# 107
C a_6293_483#0 6.4
R a_6293_483# 219
C a_5657_4411#0 8.5
R a_5657_4411# 340
C a_5777_8307#0 7.7
R a_5777_8307# 335
C a_1385_n5930#0 12.2
R a_1385_n5930# 486
C a_595_n5930#0 4.5
R a_595_n5930# 291
C a_n195_n5930#0 7.8
R a_n195_n5930# 290
C a_865_n5930#0 0.2
R a_865_n5930# 269
C a_75_n5930#0 0.0
R a_75_n5930# 269
C a_n715_n5930#0 0.0
R a_n715_n5930# 269
C a_n1505_n5930#0 2.7
R a_n1505_n5930# 974
